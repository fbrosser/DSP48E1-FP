`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:22:17 11/19/2012
// Design Name:   FPAddSub
// Module Name:   P:/FPProject/FP_AddSub/FPAddSub_tb.v
// Project Name:  FP_AddSub
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: FPAddSub
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module FPAddSub_tb;

	// Inputs
	reg clk;
	reg rst;
	reg [31:0] a;
	reg [31:0] b;
	reg operation;

	// Outputs
	wire [31:0] result;
	wire [4:0] flags;
	
	// Loop variable
	integer i;

	// Instantiate the Unit Under Test (UUT)
	FPAddSub uut (
		.clk(clk), 
		.rst(rst), 
		.a(a), 
		.b(b), 
		.operation(operation), 
		.result(result), 
		.flags(flags)
	);

	// Set up clock
	always begin
		#5 clk = ~clk;
	end

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 0;
		a = 0;
		b = 0;
		operation = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
/*
		// TEST #0
		// 8993.12 - 0.000012 = 8993
		// Expected Z = 	01000110000011001000010001111011
		#10 a = 32'b01000110000011001000010001111011; b = 32'b00110111010010010101001110011100; operation = 1'b1; $display("%b", result);

		// TEST #1
		// 8.53158062524 - 3.11224834289 = 5.41933228235
		// Expected Z = 01000000101011010110101100101100
		#10 a = 32'b01000001000010001000000101011011; b = 32'b01000000010001110010111100010100; operation = 1'b1; $display("%b", result);

		// TEST #2
		// -8.94699830093 + 2.40949324703 = -6.5375050539
		// Expected Z = 11000000110100010011001100111110
		#10 a = 32'b11000001000011110010011011101000; b = 32'b01000000000110100011010100100011; operation = 1'b0; $display("%b", result);

		// TEST #3
		// -5.82217162291 + 4.7532367122 = -1.06893491072
		// Expected Z = 10111111100010001101001011011100
		#10 a = 32'b11000000101110100100111100111011; b = 32'b01000000100110000001101010000100; operation = 1'b0; $display("%b", result);

		// TEST #4
		// 2.36803721918 - -2.82064050634 = 5.18867772552
		// Expected Z = 01000000101001100000100110100110
		#10 a = 32'b01000000000101111000110111101100; b = 32'b11000000001101001000010101100000; operation = 1'b1; $display("%b", result);

		// TEST #5
		// 3.76646645081 - 8.54622987974 = -4.77976342893
		// Expected Z = 11000000100110001111001111010010
		#10 a = 32'b01000000011100010000110111001001; b = 32'b01000001000010001011110101011100; operation = 1'b1; $display("%b", result);

		// TEST #6
		// -2.4498318859 + 5.11827801472 = 2.66844612882
		// Expected Z = 01000000001010101100011111010010
		#10 a = 32'b11000000000111001100101000001100; b = 32'b01000000101000111100100011101111; operation = 1'b0; $display("%b", result);

		// TEST #7
		// -3.2982604628 - 7.97307781549 = -11.2713382783
		// Expected Z = 11000001001101000101011101100111
		#10 a = 32'b11000000010100110001011010110011; b = 32'b01000000111111110010001101110100; operation = 1'b1; $display("%b", result);

		// TEST #8
		// 6.76606508537 + 0.854623693731 = 7.6206887791
		// Expected Z = 01000000111100111101110010101111
		#10 a = 32'b01000000110110001000001110011011; b = 32'b00111111010110101100100010011110; operation = 1'b0; $display("%b", result);

		// TEST #9
		// 9.19157019368 - -4.20144876977 = 13.3930189634
		// Expected Z = 01000001010101100100100111001110
		#10 a = 32'b01000001000100110001000010101100; b = 32'b11000000100001100111001001000101; operation = 1'b1; $display("%b", result);

		// TEST #10
		// 1.83567358255 + -8.17750207328 = -6.34182849073
		// Expected Z = 11000000110010101111000001000010
		#10 a = 32'b00111111111010101111011101011010; b = 32'b11000001000000101101011100001100; operation = 1'b0; $display("%b", result);

		for(i=0; i<=10; i=i+1) begin
			#10 $display("%b", result); 
		end 

		#100 

		#10 $finish; 
*/

// TEST #1
// 0.429198640144 + -0.702056150138 = -0.272857509994
// Expected Z = 10111110100010111011001111111011
#10 a = 32'b00111110110110111011111111101101; b = 32'b10111111001100111011100111110100; operation = 1'b0; $display("%b", result);

// TEST #2
// 0.86240205042 + -0.134426927979 = 0.727975122441
// Expected Z = 00111111001110100101110010010100
#10 a = 32'b00111111010111001100011001100001; b = 32'b10111110000010011010011100110110; operation = 1'b0; $display("%b", result);

// TEST #3
// -0.0469003428898 - 0.55705289553 = -0.60395323842
// Expected Z = 10111111000110101001110010101110
#10 a = 32'b10111101010000000001101010010011; b = 32'b00111111000011101001101100000101; operation = 1'b1; $display("%b", result);

// TEST #4
// 0.850527672867 - 0.430296703173 = 0.420230969694
// Expected Z = 00111110110101110010100010000011
#10 a = 32'b00111111010110011011110000101110; b = 32'b00111110110111000100111111011001; operation = 1'b1; $display("%b", result);

// TEST #5
// 0.846604707213 + -0.707832116689 = 0.138772590524
// Expected Z = 00111110000011100001101001100111
#10 a = 32'b00111111010110001011101100010110; b = 32'b10111111001101010011010001111100; operation = 1'b0; $display("%b", result);

// TEST #6
// 0.484029264293 + 0.382950649705 = 0.866979913998
// Expected Z = 00111111010111011111001001100101
#10 a = 32'b00111110111101111101001010101111; b = 32'b00111110110001000001001000011100; operation = 1'b0; $display("%b", result);

// TEST #7
// -0.256232203177 - 0.502954007936 = -0.759186211113
// Expected Z = 10111111010000100101101000000111
#10 a = 32'b10111110100000110011000011011110; b = 32'b00111111000000001100000110011000; operation = 1'b1; $display("%b", result);

// TEST #8
// -0.413246953076 + -0.0697155044789 = -0.482962457555
// Expected Z = 10111110111101110100011011011011
#10 a = 32'b10111110110100111001010100011011; b = 32'b10111101100011101100011100000001; operation = 1'b0; $display("%b", result);

// TEST #9
// -0.430506303883 - 0.426736061921 = -0.857242365804
// Expected Z = 10111111010110110111010000111100
#10 a = 32'b10111110110111000110101101010010; b = 32'b00111110110110100111110100100110; operation = 1'b1; $display("%b", result);

// TEST #10
// -0.731832682287 + -0.666187615042 = -1.39802029733
// Expected Z = 10111111101100101111001001010100
#10 a = 32'b10111111001110110101100101100011; b = 32'b10111111001010101000101101000110; operation = 1'b0; $display("%b", result);

// TEST #11
// -0.0603728300944 - 0.401394416206 = -0.4617672463
// Expected Z = 10111110111011000110110011000010
#10 a = 32'b10111101011101110100100110000000; b = 32'b00111110110011011000001110010010; operation = 1'b1; $display("%b", result);

// TEST #12
// -0.221730296082 + 0.251619442389 = 0.0298891463075
// Expected Z = 00111100111101001101101000010101
#10 a = 32'b10111110011000110000110101000100; b = 32'b00111110100000001101010001000011; operation = 1'b0; $display("%b", result);

// TEST #13
// -0.0938132594008 + 0.902540103395 = 0.808726843994
// Expected Z = 00111111010011110000100010111001
#10 a = 32'b10111101110000000010000100101011; b = 32'b00111111011001110000110011011110; operation = 1'b0; $display("%b", result);

// TEST #14
// 0.410328351971 + -0.602296218197 = -0.191967866226
// Expected Z = 10111110010001001001001100111001
#10 a = 32'b00111110110100100001011010001111; b = 32'b10111111000110100011000000010110; operation = 1'b0; $display("%b", result);

// TEST #15
// -0.711840021901 + -0.867110062082 = -1.57895008398
// Expected Z = 10111111110010100001101100001001
#10 a = 32'b10111111001101100011101100100110; b = 32'b10111111010111011111101011101101; operation = 1'b0; $display("%b", result);

// TEST #16
// 0.341837991461 + -0.666780954026 = -0.324942962565
// Expected Z = 10111110101001100101111011101101
#10 a = 32'b00111110101011110000010101100100; b = 32'b10111111001010101011001000101000; operation = 1'b0; $display("%b", result);

// TEST #17
// 0.701762931638 + -0.972149034859 = -0.270386103221
// Expected Z = 10111110100010100111000000001100
#10 a = 32'b00111111001100111010011010111100; b = 32'b10111111011110001101111011000010; operation = 1'b0; $display("%b", result);

// TEST #18
// -0.242543536325 - 0.607176543199 = -0.849720079525
// Expected Z = 10111111010110011000011101000001
#10 a = 32'b10111110011110000101110101010101; b = 32'b00111111000110110110111111101100; operation = 1'b1; $display("%b", result);

// TEST #19
// 0.0380149856224 + 0.347386901169 = 0.385401886792
// Expected Z = 00111110110001010101001101100101
#10 a = 32'b00111101000110111011010110011010; b = 32'b00111110101100011101110010110010; operation = 1'b0; $display("%b", result);

// TEST #20
// 0.287525296212 + -0.177245902743 = 0.110279393469
// Expected Z = 00111101111000011101101000101010
#10 a = 32'b00111110100100110011011010000100; b = 32'b10111110001101010111111111110011; operation = 1'b0; $display("%b", result);

// TEST #21
// -0.580038241506 - 0.352877820478 = -0.932916061984
// Expected Z = 10111111011011101101001110010110
#10 a = 32'b10111111000101000111110101100011; b = 32'b00111110101101001010110001100111; operation = 1'b1; $display("%b", result);

// TEST #22
// 0.597009818476 + -0.913134384131 = -0.316124565655
// Expected Z = 10111110101000011101101100010100
#10 a = 32'b00111111000110001101010110100011; b = 32'b10111111011010011100001100101101; operation = 1'b0; $display("%b", result);

// TEST #23
// -0.162184542636 + -0.208869037387 = -0.371053580023
// Expected Z = 10111110101111011111101010111100
#10 a = 32'b10111110001001100001001110110100; b = 32'b10111110010101011110000111000100; operation = 1'b0; $display("%b", result);

// TEST #24
// 0.057822270622 + 0.667497141103 = 0.725319411725
// Expected Z = 00111111001110011010111010001000
#10 a = 32'b00111101011011001101011100001100; b = 32'b00111111001010101110000100011000; operation = 1'b0; $display("%b", result);

// TEST #25
// -0.290668218956 + -0.271738722134 = -0.562406941091
// Expected Z = 10111111000011111111100111100111
#10 a = 32'b10111110100101001101001001110111; b = 32'b10111110100010110010000101010110; operation = 1'b0; $display("%b", result);

// TEST #26
// 0.596054234452 + -0.691040126065 = -0.0949858916129
// Expected Z = 10111101110000101000011111110111
#10 a = 32'b00111111000110001001011100000011; b = 32'b10111111001100001110100000000001; operation = 1'b0; $display("%b", result);

// TEST #27
// -0.329978709426 - 0.930213270191 = -1.26019197962
// Expected Z = 10111111101000010100110111111001
#10 a = 32'b10111110101010001111001011111000; b = 32'b00111111011011100010001001110101; operation = 1'b1; $display("%b", result);

// TEST #28
// -0.414966012844 + 0.700139397485 = 0.285173384641
// Expected Z = 00111110100100100000001000111111
#10 a = 32'b10111110110101000111011001101101; b = 32'b00111111001100110011110001010110; operation = 1'b0; $display("%b", result);

// TEST #29
// -0.764262575332 - -0.0686890036021 = -0.69557357173
// Expected Z = 10111111001100100001000100011100
#10 a = 32'b10111111010000111010011010110110; b = 32'b10111101100011001010110011010010; operation = 1'b1; $display("%b", result);

// TEST #30
// 0.909689647684 - -0.0443302882177 = 0.954019935902
// Expected Z = 00111111011101000011101010100111
#10 a = 32'b00111111011010001110000101101100; b = 32'b10111101001101011001001110101101; operation = 1'b1; $display("%b", result);

// TEST #31
// 0.422479032934 + -0.9675329293 = -0.545053896366
// Expected Z = 10111111000010111000100010100111
#10 a = 32'b00111110110110000100111100101100; b = 32'b10111111011101111011000000111101; operation = 1'b0; $display("%b", result);

// TEST #32
// -0.811402334357 - -0.774052341499 = -0.0373499928577
// Expected Z = 10111101000110001111110001001110
#10 a = 32'b10111111010011111011100000010000; b = 32'b10111111010001100010100001001011; operation = 1'b1; $display("%b", result);

// TEST #33
// 0.651596391088 + -0.590050606645 = 0.0615457844429
// Expected Z = 00111101011111000001011101101111
#10 a = 32'b00111111001001101100111100000101; b = 32'b10111111000101110000110110001110; operation = 1'b0; $display("%b", result);

// TEST #34
// 0.369930476848 + -0.281059091985 = 0.0888713848624
// Expected Z = 00111101101101100000001000110011
#10 a = 32'b00111110101111010110011110000111; b = 32'b10111110100011111110011011111010; operation = 1'b0; $display("%b", result);

// TEST #35
// 0.572887361768 - -0.893797361404 = 1.46668472317
// Expected Z = 00111111101110111011110001010011
#10 a = 32'b00111111000100101010100010111111; b = 32'b10111111011001001100111111100111; operation = 1'b1; $display("%b", result);

// TEST #36
// 0.358844704277 - 0.320149300468 = 0.0386954038088
// Expected Z = 00111101000111100111111100010010
#10 a = 32'b00111110101101111011101001111110; b = 32'b00111110101000111110101010011100; operation = 1'b1; $display("%b", result);

// TEST #37
// -0.640474458857 - 0.682259910111 = -1.32273436897
// Expected Z = 10111111101010010100111101011100
#10 a = 32'b10111111001000111111011000100010; b = 32'b00111111001011101010100010010110; operation = 1'b1; $display("%b", result);

// TEST #38
// 0.94466068619 + -0.708118189713 = 0.236542496477
// Expected Z = 00111110011100100011100000110010
#10 a = 32'b00111111011100011101010101001000; b = 32'b10111111001101010100011100111100; operation = 1'b0; $display("%b", result);

// TEST #39
// -0.754892127183 - 0.197302202144 = -0.952194329327
// Expected Z = 10111111011100111100001100000010
#10 a = 32'b10111111010000010100000010011100; b = 32'b00111110010010100000100110010111; operation = 1'b1; $display("%b", result);

// TEST #40
// 0.596705282497 + -0.333836897216 = 0.262868385282
// Expected Z = 00111110100001101001011010101111
#10 a = 32'b00111111000110001100000110101101; b = 32'b10111110101010101110110010101011; operation = 1'b0; $display("%b", result);

// TEST #41
// 0.863643743391 - 0.0756775715975 = 0.787966171794
// Expected Z = 00111111010010011011100000100111
#10 a = 32'b00111111010111010001011111000010; b = 32'b00111101100110101111110011011000; operation = 1'b1; $display("%b", result);

// TEST #42
// -0.224676218129 - -0.396827905098 = 0.172151686969
// Expected Z = 00111110001100000100100010001000
#10 a = 32'b10111110011001100001000110000110; b = 32'b10111110110010110010110100000111; operation = 1'b1; $display("%b", result);

// TEST #43
// 0.962138335306 - -0.868592905295 = 1.8307312406
// Expected Z = 00111111111010100101010101100111
#10 a = 32'b00111111011101100100111010110011; b = 32'b10111111010111100101110000011011; operation = 1'b1; $display("%b", result);

// TEST #44
// 0.227939519989 - 0.646227107472 = -0.418287587483
// Expected Z = 10111110110101100010100111001010
#10 a = 32'b00111110011010010110100011111010; b = 32'b00111111001001010110111100100100; operation = 1'b1; $display("%b", result);

// TEST #45
// 0.481066759666 - -0.79155932914 = 1.27262608881
// Expected Z = 00111111101000101110010101101001
#10 a = 32'b00111110111101100100111001100010; b = 32'b10111111010010101010001110100010; operation = 1'b1; $display("%b", result);

// TEST #46
// 0.225650464221 + 0.992538999942 = 1.21818946416
// Expected Z = 00111111100110111110110110100010
#10 a = 32'b00111110011001110001000011101010; b = 32'b00111111011111100001011100001001; operation = 1'b0; $display("%b", result);

// TEST #47
// 0.929324345106 + 0.166405097457 = 1.09572944256
// Expected Z = 00111111100011000100000011011101
#10 a = 32'b00111111011011011110100000110011; b = 32'b00111110001010100110011000011001; operation = 1'b0; $display("%b", result);

// TEST #48
// 0.117569447576 - -0.24376467569 = 0.361334123266
// Expected Z = 00111110101110010000000011001001
#10 a = 32'b00111101111100001100100001000000; b = 32'b10111110011110011001110101110010; operation = 1'b1; $display("%b", result);

// TEST #49
// -0.41737651817 + 0.816797127726 = 0.399420609556
// Expected Z = 00111110110011001000000011011100
#10 a = 32'b10111110110101011011001001100000; b = 32'b00111111010100010001100110011110; operation = 1'b0; $display("%b", result);

// TEST #50
// 0.739710324264 + 0.195588502991 = 0.935298827255
// Expected Z = 00111111011011110110111110111110
#10 a = 32'b00111111001111010101110110101000; b = 32'b00111110010010000100100001011010; operation = 1'b0; $display("%b", result);

// TEST #51
// 0.0923245545951 + -0.026108316574 = 0.066216238021
// Expected Z = 00111101100001111001110001100001
#10 a = 32'b00111101101111010001010010101000; b = 32'b10111100110101011110000100011100; operation = 1'b0; $display("%b", result);

// TEST #52
// 0.116034102367 - 0.935610256362 = -0.819576153995
// Expected Z = 10111111010100011100111110111110
#10 a = 32'b00111101111011011010001101001010; b = 32'b00111111011011111000010000100111; operation = 1'b1; $display("%b", result);

// TEST #53
// -0.355814414987 + 0.0537633744737 = -0.302051040514
// Expected Z = 10111110100110101010011001101111
#10 a = 32'b10111110101101100010110101001111; b = 32'b00111101010111000011011011111100; operation = 1'b0; $display("%b", result);

// TEST #54
// 0.157425693502 + 0.916109055741 = 1.07353474924
// Expected Z = 00111111100010010110100110010110
#10 a = 32'b00111110001000010011010000110011; b = 32'b00111111011010101000011000100000; operation = 1'b0; $display("%b", result);

// TEST #55
// -0.120690334958 - 0.220509108654 = -0.341199443612
// Expected Z = 10111110101011101011000110110010
#10 a = 32'b10111101111101110010110001111111; b = 32'b00111110011000011100110100100100; operation = 1'b1; $display("%b", result);

// TEST #56
// -0.00306962319164 - 0.165387622241 = -0.168457245433
// Expected Z = 10111110001011001000000000001110
#10 a = 32'b10111011010010010010101110111011; b = 32'b00111110001010010101101101011111; operation = 1'b1; $display("%b", result);

// TEST #57
// 0.456575206685 - -0.819537646902 = 1.27611285359
// Expected Z = 00111111101000110101011110101010
#10 a = 32'b00111110111010011100010000111010; b = 32'b10111111010100011100110100111000; operation = 1'b1; $display("%b", result);

// TEST #58
// 0.82231977649 - -0.820143521568 = 1.64246329806
// Expected Z = 00111111110100100011110000111101
#10 a = 32'b00111111010100101000001110001101; b = 32'b10111111010100011111010011101101; operation = 1'b1; $display("%b", result);

// TEST #59
// 0.929642827919 - -0.675869303596 = 1.60551213151
// Expected Z = 00111111110011011000000101101100
#10 a = 32'b00111111011011011111110100010011; b = 32'b10111111001011010000010111000101; operation = 1'b1; $display("%b", result);

// TEST #60
// -0.892161256724 + 0.457277296549 = -0.434883960175
// Expected Z = 10111110110111101010100100011100
#10 a = 32'b10111111011001000110010010101110; b = 32'b00111110111010100010000001000000; operation = 1'b0; $display("%b", result);

// TEST #61
// -0.446124094603 - 0.63207216232 = -1.07819625692
// Expected Z = 10111111100010100000001001010110
#10 a = 32'b10111110111001000110101001100001; b = 32'b00111111001000011100111101111011; operation = 1'b1; $display("%b", result);

// TEST #62
// 0.106070291661 - -0.181287117449 = 0.287357409111
// Expected Z = 00111110100100110010000010000011
#10 a = 32'b00111101110110010011101101100010; b = 32'b10111110001110011010001101010101; operation = 1'b1; $display("%b", result);

// TEST #63
// 0.0637573061954 + 0.992364848143 = 1.05612215434
// Expected Z = 00111111100001110010111100000011
#10 a = 32'b00111101100000101001001100110001; b = 32'b00111111011111100000101110011111; operation = 1'b0; $display("%b", result);

// TEST #64
// 0.980481367599 + -0.715634065554 = 0.264847302045
// Expected Z = 00111110100001111001101000010001
#10 a = 32'b00111111011110110000000011010100; b = 32'b10111111001101110011001111001011; operation = 1'b0; $display("%b", result);

// TEST #65
// -0.649632462323 - 0.227388576335 = -0.877021038657
// Expected Z = 10111111011000001000010001110011
#10 a = 32'b10111111001001100100111001010000; b = 32'b00111110011010001101100010001101; operation = 1'b1; $display("%b", result);

// TEST #66
// -0.00593307009037 + 0.932366697021 = 0.926433626931
// Expected Z = 00111111011011010010101011000001
#10 a = 32'b10111011110000100110101000110011; b = 32'b00111111011011101010111110010101; operation = 1'b0; $display("%b", result);

// TEST #67
// 0.256916335813 + 0.613390459801 = 0.870306795615
// Expected Z = 00111111010111101100110001101101
#10 a = 32'b00111110100000111000101010001010; b = 32'b00111111000111010000011100101000; operation = 1'b0; $display("%b", result);

// TEST #68
// 0.0327277289879 + 0.340690133113 = 0.373417862101
// Expected Z = 00111110101111110011000010100000
#10 a = 32'b00111101000001100000110110000011; b = 32'b00111110101011100110111011110000; operation = 1'b0; $display("%b", result);

// TEST #69
// 0.168860083011 - -0.899438486527 = 1.06829856954
// Expected Z = 00111111100010001011111000000010
#10 a = 32'b00111110001011001110100110101000; b = 32'b10111111011001100100000110011010; operation = 1'b1; $display("%b", result);

// TEST #70
// 0.931282967869 + -0.0329949008179 = 0.898288067051
// Expected Z = 00111111011001011111011000110101
#10 a = 32'b00111111011011100110100010010000; b = 32'b10111101000001110010010110101001; operation = 1'b0; $display("%b", result);

// TEST #71
// -0.454718601953 + -0.275245994498 = -0.729964596451
// Expected Z = 10111111001110101101111011110110
#10 a = 32'b10111110111010001101000011100000; b = 32'b10111110100011001110110100001011; operation = 1'b0; $display("%b", result);

// TEST #72
// 0.581946560041 + 0.696856224997 = 1.27880278504
// Expected Z = 00111111101000111010111111001111
#10 a = 32'b00111111000101001111101001110011; b = 32'b00111111001100100110010100101011; operation = 1'b0; $display("%b", result);

// TEST #73
// 0.35067082858 - 0.0988412463445 = 0.251829582236
// Expected Z = 00111110100000001110111111001111
#10 a = 32'b00111110101100111000101100100000; b = 32'b00111101110010100110110101001000; operation = 1'b1; $display("%b", result);

// TEST #74
// 0.859447280299 - 0.350362219106 = 0.509085061193
// Expected Z = 00111111000000100101001101100110
#10 a = 32'b00111111010111000000010010111101; b = 32'b00111110101100110110001010101101; operation = 1'b1; $display("%b", result);

// TEST #75
// -0.916190501044 + -0.632351791771 = -1.54854229281
// Expected Z = 10111111110001100011011010100010
#10 a = 32'b10111111011010101000101101110110; b = 32'b10111111001000011110000111001111; operation = 1'b0; $display("%b", result);

// TEST #76
// -0.98741953841 - -0.880172494787 = -0.107247043624
// Expected Z = 10111101110110111010010001010111
#10 a = 32'b10111111011111001100011110000111; b = 32'b10111111011000010101001011111100; operation = 1'b1; $display("%b", result);

// TEST #77
// 0.98589675274 - 0.286673469749 = 0.699223282991
// Expected Z = 00111111001100110000000001001100
#10 a = 32'b00111111011111000110001110111011; b = 32'b00111110100100101100011011011101; operation = 1'b1; $display("%b", result);

// TEST #78
// 0.412553133434 - 0.119606144597 = 0.292946988837
// Expected Z = 00111110100101011111110100100110
#10 a = 32'b00111110110100110011101000101010; b = 32'b00111101111101001111010000010001; operation = 1'b1; $display("%b", result);

// TEST #79
// -0.00360720228562 + -0.956291387738 = -0.959898590024
// Expected Z = 10111111011101011011101111101010
#10 a = 32'b10111011011011000110011011010000; b = 32'b10111111011101001100111110000011; operation = 1'b0; $display("%b", result);

// TEST #80
// -0.0365026779348 + -0.989934190012 = -1.02643686795
// Expected Z = 10111111100000110110001001001001
#10 a = 32'b10111101000101011000001111010101; b = 32'b10111111011111010110110001010100; operation = 1'b0; $display("%b", result);

// TEST #81
// -0.692307022475 + 0.128025124362 = -0.564281898113
// Expected Z = 10111111000100000111010011000111
#10 a = 32'b10111111001100010011101100001000; b = 32'b00111110000000110001100100000101; operation = 1'b0; $display("%b", result);

// TEST #82
// 0.0848902379929 - -0.0669856490082 = 0.151875887001
// Expected Z = 00111110000110111000010101011010
#10 a = 32'b00111101101011011101101011101111; b = 32'b10111101100010010010111111000110; operation = 1'b1; $display("%b", result);

// TEST #83
// -0.0447099717108 - -0.966960317468 = 0.922250345758
// Expected Z = 00111111011011000001100010011001
#10 a = 32'b10111101001101110010000111001110; b = 32'b10111111011101111000101010110110; operation = 1'b1; $display("%b", result);

// TEST #84
// 0.0301132211612 + 0.727532638712 = 0.757645859873
// Expected Z = 00111111010000011111010100010100
#10 a = 32'b00111100111101101011000000000001; b = 32'b00111111001110100011111110010100; operation = 1'b0; $display("%b", result);

// TEST #85
// 0.215582516895 - -0.754395444081 = 0.969977960976
// Expected Z = 00111111011110000101000001111010
#10 a = 32'b00111110010111001100000110101010; b = 32'b10111111010000010010000000001111; operation = 1'b1; $display("%b", result);

// TEST #86
// 0.68934133774 + 0.764717710714 = 1.45405904845
// Expected Z = 00111111101110100001111010011011
#10 a = 32'b00111111001100000111100010101101; b = 32'b00111111010000111100010010001010; operation = 1'b0; $display("%b", result);

// TEST #87
// -0.845917898482 - 0.803557943179 = -1.64947584166
// Expected Z = 10111111110100110010001000000110
#10 a = 32'b10111111010110001000111000010011; b = 32'b00111111010011011011010111111001; operation = 1'b1; $display("%b", result);

// TEST #88
// -0.463261738595 - 0.181907995083 = -0.645169733678
// Expected Z = 10111111001001010010100111011000
#10 a = 32'b10111110111011010011000010100101; b = 32'b00111110001110100100011000010111; operation = 1'b1; $display("%b", result);

// TEST #89
// 0.425192395955 + -0.0191897401051 = 0.40600265585
// Expected Z = 00111110110011111101111110010101
#10 a = 32'b00111110110110011011001011010001; b = 32'b10111100100111010011001111001101; operation = 1'b0; $display("%b", result);

// TEST #90
// -0.134183677929 - -0.476269609408 = 0.342085931478
// Expected Z = 00111110101011110010010111100011
#10 a = 32'b10111110000010010110011101110010; b = 32'b10111110111100111101100110011100; operation = 1'b1; $display("%b", result);

// TEST #91
// -0.4184062307 - 0.468968027021 = -0.887374257721
// Expected Z = 10111111011000110010101011110110
#10 a = 32'b10111110110101100011100101010111; b = 32'b00111110111100000001110010010100; operation = 1'b1; $display("%b", result);

// TEST #92
// 0.73299904045 + -0.983440282839 = -0.250441242389
// Expected Z = 10111110100000000011100111010110
#10 a = 32'b00111111001110111010010111010011; b = 32'b10111111011110111100001010111110; operation = 1'b0; $display("%b", result);

// TEST #93
// 0.841236740299 - -0.55445543143 = 1.39569217173
// Expected Z = 00111111101100101010011000001011
#10 a = 32'b00111111010101110101101101001010; b = 32'b10111111000011011111000011001011; operation = 1'b1; $display("%b", result);

// TEST #94
// -0.664660427235 + -0.824865307038 = -1.48952573427
// Expected Z = 10111111101111101010100011000111
#10 a = 32'b10111111001010100010011100110000; b = 32'b10111111010100110010101001011111; operation = 1'b0; $display("%b", result);

// TEST #95
// 0.946861077128 + -0.389836095299 = 0.557024981829
// Expected Z = 00111111000011101001100100110000
#10 a = 32'b00111111011100100110010101111101; b = 32'b10111110110001111001100010011001; operation = 1'b0; $display("%b", result);

// TEST #96
// 0.613950173428 - 0.880552558225 = -0.266602384797
// Expected Z = 10111110100010001000000000011100
#10 a = 32'b00111111000111010010101111010111; b = 32'b00111111011000010110101111100100; operation = 1'b1; $display("%b", result);

// TEST #97
// -0.970523377289 - 0.475259142416 = -1.4457825197
// Expected Z = 10111111101110010000111101100111
#10 a = 32'b10111111011110000111010000111000; b = 32'b00111110111100110101010100101011; operation = 1'b1; $display("%b", result);

// TEST #98
// -0.202255406072 + 0.900902324206 = 0.698646918134
// Expected Z = 00111111001100101101101010000110
#10 a = 32'b10111110010011110001110000001011; b = 32'b00111111011001101010000110001001; operation = 1'b0; $display("%b", result);

// TEST #99
// -0.139698244324 - -0.73315448882 = 0.593456244496
// Expected Z = 00111111000101111110110011000000
#10 a = 32'b10111110000011110000110100001110; b = 32'b10111111001110111011000000000011; operation = 1'b1; $display("%b", result);

// TEST #100
// 0.230589714643 + 0.375276307349 = 0.605866021992
// Expected Z = 00111111000110110001101000001001
#10 a = 32'b00111110011011000001111110110110; b = 32'b00111110110000000010010000110111; operation = 1'b0; $display("%b", result);

// TEST #101
// 519.065976251 + 288.579844274 = 807.645820524
// Expected Z = 01000100010010011110100101010101
#10 a = 32'b01000100000000011100010000111001; b = 32'b01000011100100000100101000111000; operation = 1'b0; $display("%b", result);

// TEST #102
// -336.600984741 - -533.162049286 = 196.561064545
// Expected Z = 01000011010001001000111110100010
#10 a = 32'b11000011101010000100110011101101; b = 32'b11000100000001010100101001011111; operation = 1'b1; $display("%b", result);

// TEST #103
// -672.351676402 + 353.78488429 = -318.566792112
// Expected Z = 11000011100111110100100010001101
#10 a = 32'b11000100001010000001011010000010; b = 32'b01000011101100001110010001110111; operation = 1'b0; $display("%b", result);

// TEST #104
// 336.481199551 - -778.298764773 = 1114.77996432
// Expected Z = 01000100100010110101100011110101
#10 a = 32'b01000011101010000011110110011000; b = 32'b11000100010000101001001100011111; operation = 1'b1; $display("%b", result);

// TEST #105
// -639.866452142 + -124.012511399 = -763.878963541
// Expected Z = 11000100001111101111100001000001
#10 a = 32'b11000100000111111111011101110100; b = 32'b11000010111110000000011001101000; operation = 1'b0; $display("%b", result);

// TEST #106
// -924.097534917 - 346.830316789 = -1270.92785171
// Expected Z = 11000100100111101101110110110001
#10 a = 32'b11000100011001110000011000111110; b = 32'b01000011101011010110101001001000; operation = 1'b1; $display("%b", result);

// TEST #107
// 898.655580954 - 259.280915137 = 639.374665817
// Expected Z = 01000100000111111101011111111011
#10 a = 32'b01000100011000001010100111110101; b = 32'b01000011100000011010001111110101; operation = 1'b1; $display("%b", result);

// TEST #108
// -551.827110181 - 993.478020955 = -1545.30513114
// Expected Z = 11000100110000010010100111000100
#10 a = 32'b11000100000010011111010011101111; b = 32'b01000100011110000101111010011000; operation = 1'b1; $display("%b", result);

// TEST #109
// -969.724984397 - -766.261846138 = -203.463138259
// Expected Z = 11000011010010110111011010010000
#10 a = 32'b11000100011100100110111001100110; b = 32'b11000100001111111001000011000010; operation = 1'b1; $display("%b", result);

// TEST #110
// 768.859749617 + 534.057774659 = 1302.91752428
// Expected Z = 01000100101000101101110101011100
#10 a = 32'b01000100010000000011011100000110; b = 32'b01000100000001011000001110110011; operation = 1'b0; $display("%b", result);

// TEST #111
// 290.654999761 + -496.070824055 = -205.415824294
// Expected Z = 11000011010011010110101001110011
#10 a = 32'b01000011100100010101001111010111; b = 32'b11000011111110000000100100010001; operation = 1'b0; $display("%b", result);

// TEST #112
// -288.999917906 + 463.36538673 = 174.365468824
// Expected Z = 01000011001011100101110110001111
#10 a = 32'b11000011100100000111111111111101; b = 32'b01000011111001111010111011000101; operation = 1'b0; $display("%b", result);

// TEST #113
// 699.556738626 - 155.781758099 = 543.774980527
// Expected Z = 01000100000001111111000110011001
#10 a = 32'b01000100001011101110001110100010; b = 32'b01000011000110111100100000100001; operation = 1'b1; $display("%b", result);

// TEST #114
// 44.4148565778 - 916.197159576 = -871.782302999
// Expected Z = 11000100010110011111001000010001
#10 a = 32'b01000010001100011010100011010000; b = 32'b01000100011001010000110010011110; operation = 1'b1; $display("%b", result);

// TEST #115
// -799.799107267 - -344.966836681 = -454.832270585
// Expected Z = 11000011111000110110101010001000
#10 a = 32'b11000100010001111111001100100101; b = 32'b11000011101011000111101111000001; operation = 1'b1; $display("%b", result);

// TEST #116
// 368.070563925 + -832.04690753 = -463.976343605
// Expected Z = 11000011111001111111110011111001
#10 a = 32'b01000011101110000000100100001000; b = 32'b11000100010100000000001100000001; operation = 1'b0; $display("%b", result);

// TEST #117
// 267.426779756 + -129.800003882 = 137.626775874
// Expected Z = 01000011000010011010000001110100
#10 a = 32'b01000011100001011011011010100001; b = 32'b11000011000000011100110011001101; operation = 1'b0; $display("%b", result);

// TEST #118
// 674.4165915 + -537.232338644 = 137.184252856
// Expected Z = 01000011000010010010111100101011
#10 a = 32'b01000100001010001001101010101001; b = 32'b11000100000001100100111011011111; operation = 1'b0; $display("%b", result);

// TEST #119
// 127.986308217 - -209.398417253 = 337.38472547
// Expected Z = 01000011101010001011000100111111
#10 a = 32'b01000010111111111111100011111101; b = 32'b11000011010100010110010111111111; operation = 1'b1; $display("%b", result);

// TEST #120
// -227.088717625 - 743.971054955 = -971.059772581
// Expected Z = 11000100011100101100001111010011
#10 a = 32'b11000011011000110001011010110110; b = 32'b01000100001110011111111000100110; operation = 1'b1; $display("%b", result);

// TEST #121
// 488.394212637 + -586.89674732 = -98.5025346832
// Expected Z = 11000010110001010000000101001100
#10 a = 32'b01000011111101000011001001110110; b = 32'b11000100000100101011100101100100; operation = 1'b0; $display("%b", result);

// TEST #122
// 35.6145739953 + 877.091628421 = 912.706202416
// Expected Z = 01000100011001000010110100110010
#10 a = 32'b01000010000011100111010101010011; b = 32'b01000100010110110100010111011101; operation = 1'b0; $display("%b", result);

// TEST #123
// 624.905240183 - 181.489977796 = 443.415262387
// Expected Z = 01000011110111011011010100100111
#10 a = 32'b01000100000111000011100111101111; b = 32'b01000011001101010111110101101111; operation = 1'b1; $display("%b", result);

// TEST #124
// 917.623780078 - -673.835932491 = 1591.45971257
// Expected Z = 01000100110001101110111010110110
#10 a = 32'b01000100011001010110011111101100; b = 32'b11000100001010000111010110000000; operation = 1'b1; $display("%b", result);

// TEST #125
// 570.410844977 - 867.395120949 = -296.984275973
// Expected Z = 11000011100101000111110111111101
#10 a = 32'b01000100000011101001101001001011; b = 32'b01000100010110001101100101001010; operation = 1'b1; $display("%b", result);

// TEST #126
// -867.415039605 - 928.080070876 = -1795.49511048
// Expected Z = 11000100111000000110111111011000
#10 a = 32'b11000100010110001101101010010000; b = 32'b01000100011010000000010100100000; operation = 1'b1; $display("%b", result);

// TEST #127
// -398.389155086 + -502.941985463 = -901.331140549
// Expected Z = 11000100011000010101010100110001
#10 a = 32'b11000011110001110011000111010000; b = 32'b11000011111110110111100010010011; operation = 1'b0; $display("%b", result);

// TEST #128
// 248.871326619 - 194.64323519 = 54.2280914287
// Expected Z = 01000010010110001110100110010001
#10 a = 32'b01000011011110001101111100001111; b = 32'b01000011010000101010010010101011; operation = 1'b1; $display("%b", result);

// TEST #129
// 289.67153102 - -149.845778345 = 439.517309364
// Expected Z = 01000011110110111100001000110111
#10 a = 32'b01000011100100001101010111110101; b = 32'b11000011000101011101100010000101; operation = 1'b1; $display("%b", result);

// TEST #130
// -484.280379618 + -733.752135999 = -1218.03251562
// Expected Z = 11000100100110000100000100001010
#10 a = 32'b11000011111100100010001111100011; b = 32'b11000100001101110111000000100011; operation = 1'b0; $display("%b", result);

// TEST #131
// 973.801738861 - 902.482883787 = 71.3188550743
// Expected Z = 01000010100011101010001101000001
#10 a = 32'b01000100011100110111001101010000; b = 32'b01000100011000011001111011101000; operation = 1'b1; $display("%b", result);

// TEST #132
// -91.6746012426 - -222.304516372 = 130.629915129
// Expected Z = 01000011000000101010000101000010
#10 a = 32'b11000010101101110101100101100101; b = 32'b11000011010111100100110111110101; operation = 1'b1; $display("%b", result);

// TEST #133
// -230.890794795 + -293.598215167 = -524.489009962
// Expected Z = 11000100000000110001111101001100
#10 a = 32'b11000011011001101110010000001011; b = 32'b11000011100100101100110010010010; operation = 1'b0; $display("%b", result);

// TEST #134
// 450.893546159 - -656.9826282 = 1107.87617436
// Expected Z = 01000100100010100111110000001010
#10 a = 32'b01000011111000010111001001100000; b = 32'b11000100001001000011111011100011; operation = 1'b1; $display("%b", result);

// TEST #135
// 847.945374185 - 95.9759204574 = 751.969453728
// Expected Z = 01000100001110111111111000001100
#10 a = 32'b01000100010100111111110010000001; b = 32'b01000010101111111111001110101100; operation = 1'b1; $display("%b", result);

// TEST #136
// 733.785261487 + 722.659868429 = 1456.44512992
// Expected Z = 01000100101101100000111000111111
#10 a = 32'b01000100001101110111001001000010; b = 32'b01000100001101001010101000111011; operation = 1'b0; $display("%b", result);

// TEST #137
// 586.622398384 + 302.372737231 = 888.995135615
// Expected Z = 01000100010111100011111110110000
#10 a = 32'b01000100000100101010011111010101; b = 32'b01000011100101110010111110110110; operation = 1'b0; $display("%b", result);

// TEST #138
// 843.875523161 - 206.540499194 = 637.335023967
// Expected Z = 01000100000111110101010101110001
#10 a = 32'b01000100010100101111100000001001; b = 32'b01000011010011101000101001011110; operation = 1'b1; $display("%b", result);

// TEST #139
// -275.913145561 + 406.073230774 = 130.160085213
// Expected Z = 01000011000000100010100011111011
#10 a = 32'b11000011100010011111010011100010; b = 32'b01000011110010110000100101100000; operation = 1'b0; $display("%b", result);

// TEST #140
// -374.827846813 + 951.965869357 = 577.138022544
// Expected Z = 01000100000100000100100011010101
#10 a = 32'b11000011101110110110100111110111; b = 32'b01000100011011011111110111010001; operation = 1'b0; $display("%b", result);

// TEST #141
// -330.990451383 - -632.144155795 = 301.153704412
// Expected Z = 01000011100101101001001110101101
#10 a = 32'b11000011101001010111111011000111; b = 32'b11000100000111100000100100111010; operation = 1'b1; $display("%b", result);

// TEST #142
// 165.000040976 - 365.282464654 = -200.282423678
// Expected Z = 11000011010010000100100001001101
#10 a = 32'b01000011001001010000000000000011; b = 32'b01000011101101101010010000101000; operation = 1'b1; $display("%b", result);

// TEST #143
// -843.257434535 - 475.037259015 = -1318.29469355
// Expected Z = 11000100101001001100100101101110
#10 a = 32'b11000100010100101101000001111010; b = 32'b01000011111011011000010011000101; operation = 1'b1; $display("%b", result);

// TEST #144
// -921.603800123 + -412.740974874 = -1334.344775
// Expected Z = 11000100101001101100101100001000
#10 a = 32'b11000100011001100110011010100101; b = 32'b11000011110011100101111011011000; operation = 1'b0; $display("%b", result);

// TEST #145
// -26.9775904001 + -220.809717252 = -247.787307652
// Expected Z = 11000011011101111100100110001101
#10 a = 32'b11000001110101111101001000011011; b = 32'b11000011010111001100111101001010; operation = 1'b0; $display("%b", result);

// TEST #146
// -643.817521579 + 244.216259222 = -399.601262357
// Expected Z = 11000011110001111100110011110110
#10 a = 32'b11000100001000001111010001010010; b = 32'b01000011011101000011011101011101; operation = 1'b0; $display("%b", result);

// TEST #147
// 660.933748473 + -711.262236614 = -50.3284881418
// Expected Z = 11000010010010010101000001011111
#10 a = 32'b01000100001001010011101111000011; b = 32'b11000100001100011101000011001000; operation = 1'b0; $display("%b", result);

// TEST #148
// -499.526046889 + -915.847046804 = -1415.37309369
// Expected Z = 11000100101100001110101111110000
#10 a = 32'b11000011111110011100001101010110; b = 32'b11000100011001001111011000110110; operation = 1'b0; $display("%b", result);

// TEST #149
// 722.586796422 - 551.697888362 = 170.888908061
// Expected Z = 01000011001010101110001110001111
#10 a = 32'b01000100001101001010010110001110; b = 32'b01000100000010011110110010101010; operation = 1'b1; $display("%b", result);

// TEST #150
// 613.151399025 - 394.875524111 = 218.275874914
// Expected Z = 01000011010110100100011010100000
#10 a = 32'b01000100000110010100100110110001; b = 32'b01000011110001010111000000010001; operation = 1'b1; $display("%b", result);

// TEST #151
// -851.194011513 + -54.6099938532 = -905.804005367
// Expected Z = 11000100011000100111001101110101
#10 a = 32'b11000100010101001100110001101011; b = 32'b11000010010110100111000010100010; operation = 1'b0; $display("%b", result);

// TEST #152
// 725.061688253 + 866.443798377 = 1591.50548663
// Expected Z = 01000100110001101111000000101101
#10 a = 32'b01000100001101010100001111110011; b = 32'b01000100010110001001110001100111; operation = 1'b0; $display("%b", result);

// TEST #153
// 968.782967243 + 999.5997369 = 1968.38270414
// Expected Z = 01000100111101100000110000111111
#10 a = 32'b01000100011100100011001000011100; b = 32'b01000100011110011110011001100010; operation = 1'b0; $display("%b", result);

// TEST #154
// 377.425858375 + -436.927172495 = -59.5013141198
// Expected Z = 11000010011011100000000101011000
#10 a = 32'b01000011101111001011011010000011; b = 32'b11000011110110100111011010101110; operation = 1'b0; $display("%b", result);

// TEST #155
// -393.476038241 - 135.623693575 = -529.099731816
// Expected Z = 11000100000001000100011001100010
#10 a = 32'b11000011110001001011110011101111; b = 32'b01000011000001111001111110101010; operation = 1'b1; $display("%b", result);

// TEST #156
// -291.467771472 - 430.061709369 = -721.529480841
// Expected Z = 11000100001101000110000111100011
#10 a = 32'b11000011100100011011101111100000; b = 32'b01000011110101110000011111100110; operation = 1'b1; $display("%b", result);

// TEST #157
// -13.5716254095 + -243.901387486 = -257.473012896
// Expected Z = 11000011100000001011110010001100
#10 a = 32'b11000001010110010010010101100001; b = 32'b11000011011100111110011011000001; operation = 1'b0; $display("%b", result);

// TEST #158
// -392.557012591 - -328.755854049 = -63.8011585416
// Expected Z = 11000010011111110011010001100011
#10 a = 32'b11000011110001000100011101001100; b = 32'b11000011101001000110000011000000; operation = 1'b1; $display("%b", result);

// TEST #159
// -620.988263889 + -937.954484329 = -1558.94274822
// Expected Z = 11000100110000101101111000101011
#10 a = 32'b11000100000110110011111101000000; b = 32'b11000100011010100111110100010110; operation = 1'b0; $display("%b", result);

// TEST #160
// 728.048686658 + -20.8612342022 = 707.187452455
// Expected Z = 01000100001100001100101111111111
#10 a = 32'b01000100001101100000001100011110; b = 32'b11000001101001101110001111001111; operation = 1'b0; $display("%b", result);

// TEST #161
// -649.579542129 + 795.029927091 = 145.450384962
// Expected Z = 01000011000100010111001101001100
#10 a = 32'b11000100001000100110010100010111; b = 32'b01000100010001101100000111101010; operation = 1'b0; $display("%b", result);

// TEST #162
// -613.490079505 - -122.709590863 = -490.780488642
// Expected Z = 11000011111101010110001111100111
#10 a = 32'b11000100000110010101111101011101; b = 32'b11000010111101010110101101001111; operation = 1'b1; $display("%b", result);

// TEST #163
// 370.004149312 - -576.593203711 = 946.597353024
// Expected Z = 01000100011011001010011000111011
#10 a = 32'b01000011101110010000000010001000; b = 32'b11000100000100000010010111110111; operation = 1'b1; $display("%b", result);

// TEST #164
// -897.22697561 + 940.821902531 = 43.5949269214
// Expected Z = 01000010001011100110000100110101
#10 a = 32'b11000100011000000100111010000111; b = 32'b01000100011010110011010010011010; operation = 1'b0; $display("%b", result);

// TEST #165
// -755.219464591 - 266.058981293 = -1021.27844588
// Expected Z = 11000100011111110101000111010010
#10 a = 32'b11000100001111001100111000001100; b = 32'b01000011100001010000011110001101; operation = 1'b1; $display("%b", result);

// TEST #166
// -565.500801756 - -614.965736279 = 49.4649345236
// Expected Z = 01000010010001011101110000011000
#10 a = 32'b11000100000011010110000000001101; b = 32'b11000100000110011011110111001111; operation = 1'b1; $display("%b", result);

// TEST #167
// 878.514366013 + -476.685154049 = 401.829211964
// Expected Z = 01000011110010001110101000100100
#10 a = 32'b01000100010110111010000011101011; b = 32'b11000011111011100101011110110011; operation = 1'b0; $display("%b", result);

// TEST #168
// -51.8475701854 - 52.236548128 = -104.084118313
// Expected Z = 11000010110100000010101100010010
#10 a = 32'b11000010010011110110001111101001; b = 32'b01000010010100001111001000111010; operation = 1'b1; $display("%b", result);

// TEST #169
// 656.807998824 + -20.2038458185 = 636.604153006
// Expected Z = 01000100000111110010011010101010
#10 a = 32'b01000100001001000011001110110110; b = 32'b11000001101000011010000101111010; operation = 1'b0; $display("%b", result);

// TEST #170
// 186.886093267 - 447.278009414 = -260.391916146
// Expected Z = 11000011100000100011001000101010
#10 a = 32'b01000011001110101110001011010111; b = 32'b01000011110111111010001110010110; operation = 1'b1; $display("%b", result);

// TEST #171
// 488.007528238 + -574.395660469 = -86.3881322309
// Expected Z = 11000010101011001100011010111001
#10 a = 32'b01000011111101000000000011110111; b = 32'b11000100000011111001100101010011; operation = 1'b0; $display("%b", result);

// TEST #172
// -626.0766235 + 552.280464889 = -73.7961586103
// Expected Z = 11000010100100111001011110100010
#10 a = 32'b11000100000111001000010011100111; b = 32'b01000100000010100001000111110011; operation = 1'b0; $display("%b", result);

// TEST #173
// -723.83458639 - 449.140927997 = -1172.97551439
// Expected Z = 11000100100100101001111100110111
#10 a = 32'b11000100001101001111010101101010; b = 32'b01000011111000001001001000001010; operation = 1'b1; $display("%b", result);

// TEST #174
// -488.815452338 + 643.912849196 = 155.097396858
// Expected Z = 01000011000110110001100011101111
#10 a = 32'b11000011111101000110100001100001; b = 32'b01000100001000001111101001101100; operation = 1'b0; $display("%b", result);

// TEST #175
// 991.448057799 - -291.529991291 = 1282.97804909
// Expected Z = 01000100101000000101111101001100
#10 a = 32'b01000100011101111101110010101101; b = 32'b11000011100100011100001111010111; operation = 1'b1; $display("%b", result);

// TEST #176
// 51.1795887906 - -79.9157819301 = 131.095370721
// Expected Z = 01000011000000110001100001101010
#10 a = 32'b01000010010011001011011111100110; b = 32'b11000010100111111101010011100001; operation = 1'b1; $display("%b", result);

// TEST #177
// 305.385899351 + -976.323838345 = -670.937938994
// Expected Z = 11000100001001111011110000000111
#10 a = 32'b01000011100110001011000101100101; b = 32'b11000100011101000001010010111010; operation = 1'b0; $display("%b", result);

// TEST #178
// -375.44557135 + -696.551689237 = -1071.99726059
// Expected Z = 11000100100001011111111111101010
#10 a = 32'b11000011101110111011100100001000; b = 32'b11000100001011100010001101001111; operation = 1'b0; $display("%b", result);

// TEST #179
// -287.878595504 + 146.341102011 = -141.537493493
// Expected Z = 11000011000011011000100110011001
#10 a = 32'b11000011100011111111000001110110; b = 32'b01000011000100100101011101010010; operation = 1'b0; $display("%b", result);

// TEST #180
// 109.300594428 - 596.517038138 = -487.216443709
// Expected Z = 11000011111100111001101110110100
#10 a = 32'b01000010110110101001100111101000; b = 32'b01000100000101010010000100010111; operation = 1'b1; $display("%b", result);

// TEST #181
// 56.9393437991 + -863.398397202 = -806.459053403
// Expected Z = 11000100010010011001110101100001
#10 a = 32'b01000010011000111100000111100011; b = 32'b11000100010101111101100101111111; operation = 1'b0; $display("%b", result);

// TEST #182
// -328.980106695 - -663.959767545 = 334.97966085
// Expected Z = 01000011101001110111110101100110
#10 a = 32'b11000011101001000111110101110100; b = 32'b11000100001001011111110101101101; operation = 1'b1; $display("%b", result);

// TEST #183
// -162.884609722 + -241.18098352 = -404.065593242
// Expected Z = 11000011110010100000100001100101
#10 a = 32'b11000011001000101110001001110110; b = 32'b11000011011100010010111001010101; operation = 1'b0; $display("%b", result);

// TEST #184
// 359.290791326 + -906.633032112 = -547.342240786
// Expected Z = 11000100000010001101010111100111
#10 a = 32'b01000011101100111010010100111001; b = 32'b11000100011000101010100010000100; operation = 1'b0; $display("%b", result);

// TEST #185
// 826.879133584 + -571.270050862 = 255.609082722
// Expected Z = 01000011011111111001101111101101
#10 a = 32'b01000100010011101011100001000100; b = 32'b11000100000011101101000101001001; operation = 1'b0; $display("%b", result);

// TEST #186
// -838.947457808 - 824.768356288 = -1663.7158141
// Expected Z = 11000100110011111111011011101000
#10 a = 32'b11000100010100011011110010100011; b = 32'b01000100010011100011000100101101; operation = 1'b1; $display("%b", result);

// TEST #187
// 711.825124651 - 255.09526508 = 456.729859571
// Expected Z = 01000011111001000101110101101100
#10 a = 32'b01000100001100011111010011001111; b = 32'b01000011011111110001100001100011; operation = 1'b1; $display("%b", result);

// TEST #188
// 543.930983222 + 256.070829554 = 800.001812776
// Expected Z = 01000100010010000000000000011110
#10 a = 32'b01000100000001111111101110010101; b = 32'b01000011100000000000100100010001; operation = 1'b0; $display("%b", result);

// TEST #189
// -948.387969854 + -197.197847252 = -1145.58581711
// Expected Z = 11000100100011110011001010111111
#10 a = 32'b11000100011011010001100011010100; b = 32'b11000011010001010011001010100110; operation = 1'b0; $display("%b", result);

// TEST #190
// -575.492048569 - -197.844417491 = -377.647631078
// Expected Z = 11000011101111001101001011100110
#10 a = 32'b11000100000011111101111101111110; b = 32'b11000011010001011101100000101100; operation = 1'b1; $display("%b", result);

// TEST #191
// 39.6238845048 + -659.791759284 = -620.167874779
// Expected Z = 11000100000110110000101010111110
#10 a = 32'b01000010000111100111111011011100; b = 32'b11000100001001001111001010101100; operation = 1'b0; $display("%b", result);

// TEST #192
// -362.805746664 - 84.127650008 = -446.933396672
// Expected Z = 11000011110111110111011101111010
#10 a = 32'b11000011101101010110011100100011; b = 32'b01000010101010000100000101011011; operation = 1'b1; $display("%b", result);

// TEST #193
// 129.315280966 - -994.330898288 = 1123.64617925
// Expected Z = 01000100100011000111010010101110
#10 a = 32'b01000011000000010101000010110110; b = 32'b11000100011110001001010100101101; operation = 1'b1; $display("%b", result);

// TEST #194
// 137.629929035 + -376.690288823 = -239.060359788
// Expected Z = 11000011011011110000111101110100
#10 a = 32'b01000011000010011010000101000011; b = 32'b11000011101111000101100001011011; operation = 1'b0; $display("%b", result);

// TEST #195
// 468.804722378 + 960.764937911 = 1429.56966029
// Expected Z = 01000100101100101011001000111011
#10 a = 32'b01000011111010100110011100000001; b = 32'b01000100011100000011000011110101; operation = 1'b0; $display("%b", result);

// TEST #196
// -442.732441556 - -563.334044335 = 120.601602778
// Expected Z = 01000010111100010011010000000101
#10 a = 32'b11000011110111010101110111000001; b = 32'b11000100000011001101010101100001; operation = 1'b1; $display("%b", result);

// TEST #197
// -892.344264245 - -161.212968552 = -731.131295694
// Expected Z = 11000100001101101100100001100111
#10 a = 32'b11000100010111110001011000001000; b = 32'b11000011001000010011011010000101; operation = 1'b1; $display("%b", result);

// TEST #198
// 532.250046974 + -448.586782524 = 83.6632644496
// Expected Z = 01000010101001110101001110010111
#10 a = 32'b01000100000001010001000000000001; b = 32'b11000011111000000100101100011100; operation = 1'b0; $display("%b", result);

// TEST #199
// 530.930756985 - -181.989520774 = 712.920277759
// Expected Z = 01000100001100100011101011100110
#10 a = 32'b01000100000001001011101110010010; b = 32'b11000011001101011111110101010001; operation = 1'b1; $display("%b", result);

// TEST #200
// 128.048594794 - -732.756474226 = 860.80506902
// Expected Z = 01000100010101110011001110000110
#10 a = 32'b01000011000000000000110001110001; b = 32'b11000100001101110011000001101010; operation = 1'b1; $display("%b", result);

// TEST #201
// 0.987064259885 + -112.178973928 = -111.191909668
// Expected Z = 11000010110111100110001001000010
#10 a = 32'b00111111011111001011000000111110; b = 32'b11000010111000000101101110100010; operation = 1'b0; $display("%b", result);

// TEST #202
// -0.26423463325 - -685.878022055 = 685.613787422
// Expected Z = 01000100001010110110011101001000
#10 a = 32'b10111110100001110100100111000011; b = 32'b11000100001010110111100000110010; operation = 1'b1; $display("%b", result);

// TEST #203
// -0.39357684383 - -381.649936015 = 381.256359171
// Expected Z = 01000011101111101010000011010000
#10 a = 32'b10111110110010011000001011100111; b = 32'b11000011101111101101001100110001; operation = 1'b1; $display("%b", result);

// TEST #204
// -0.146099548663 + -240.714004995 = -240.860104544
// Expected Z = 11000011011100001101110000110000
#10 a = 32'b10111110000101011001101100011111; b = 32'b11000011011100001011011011001001; operation = 1'b0; $display("%b", result);

// TEST #205
// -0.541659573373 - -286.239929454 = 285.698269881
// Expected Z = 01000011100011101101100101100001
#10 a = 32'b10111111000010101010101000110100; b = 32'b11000011100011110001111010110110; operation = 1'b1; $display("%b", result);

// TEST #206
// 0.826332088967 - 825.159819002 = -824.333486913
// Expected Z = 11000100010011100001010101011000
#10 a = 32'b00111111010100111000101010000000; b = 32'b01000100010011100100101000111010; operation = 1'b1; $display("%b", result);

// TEST #207
// -0.925182400532 - 569.781835782 = -570.707018182
// Expected Z = 11000100000011101010110101000000
#10 a = 32'b10111111011011001101100011000001; b = 32'b01000100000011100111001000001010; operation = 1'b1; $display("%b", result);

// TEST #208
// 0.804638437553 - -582.023830084 = 582.828468522
// Expected Z = 01000100000100011011010100000110
#10 a = 32'b00111111010011011111110011001001; b = 32'b11000100000100011000000110000110; operation = 1'b1; $display("%b", result);

// TEST #209
// 0.201346878512 - -495.687737117 = 495.889083996
// Expected Z = 01000011111101111111000111001110
#10 a = 32'b00111110010011100010110111100000; b = 32'b11000011111101111101100000001000; operation = 1'b1; $display("%b", result);

// TEST #210
// -0.987863546602 + 357.053568857 = 356.065705311
// Expected Z = 01000011101100100000100001101001
#10 a = 32'b10111111011111001110010010100000; b = 32'b01000011101100101000011011011011; operation = 1'b0; $display("%b", result);

// TEST #211
// -0.516105977341 - -879.291762234 = 878.775656257
// Expected Z = 01000100010110111011000110100100
#10 a = 32'b10111111000001000001111110000101; b = 32'b11000100010110111101001010101100; operation = 1'b1; $display("%b", result);

// TEST #212
// -0.0890908344861 - -75.9188787119 = 75.8297878774
// Expected Z = 01000010100101111010100011011010
#10 a = 32'b10111101101101100111010101000001; b = 32'b11000010100101111101011001110111; operation = 1'b1; $display("%b", result);

// TEST #213
// 0.203033955437 - 827.718708223 = -827.515674268
// Expected Z = 11000100010011101110000100000001
#10 a = 32'b00111110010011111110100000100010; b = 32'b01000100010011101110110111111111; operation = 1'b1; $display("%b", result);

// TEST #214
// 0.946123144459 - -386.400984396 = 387.34710754
// Expected Z = 01000011110000011010110001101110
#10 a = 32'b00111111011100100011010100100000; b = 32'b11000011110000010011001101010011; operation = 1'b1; $display("%b", result);

// TEST #215
// -0.957332785185 + 152.646851626 = 151.689518841
// Expected Z = 01000011000101111011000010000100
#10 a = 32'b10111111011101010001001111000011; b = 32'b01000011000110001010010110011000; operation = 1'b0; $display("%b", result);

// TEST #216
// 0.0418448172949 + -423.427816208 = -423.385971391
// Expected Z = 11000011110100111011000101101000
#10 a = 32'b00111101001010110110010101111001; b = 32'b11000011110100111011011011000011; operation = 1'b0; $display("%b", result);

// TEST #217
// 0.412895376165 - 626.163549291 = -625.750653915
// Expected Z = 11000100000111000111000000001011
#10 a = 32'b00111110110100110110011100000110; b = 32'b01000100000111001000101001111000; operation = 1'b1; $display("%b", result);

// TEST #218
// 0.0339284117145 - 767.838351554 = -767.804423142
// Expected Z = 11000100001111111111001101111100
#10 a = 32'b00111101000010101111100010000101; b = 32'b01000100001111111111010110101000; operation = 1'b1; $display("%b", result);

// TEST #219
// -0.846718849143 + 177.74619192 = 176.89947307
// Expected Z = 01000011001100001110011001000100
#10 a = 32'b10111111010110001100001010010001; b = 32'b01000011001100011011111100000110; operation = 1'b0; $display("%b", result);

// TEST #220
// -0.355337153716 - -16.2216351581 = 15.8662980044
// Expected Z = 01000001011111011101110001011011
#10 a = 32'b10111110101101011110111011000000; b = 32'b11000001100000011100010111101001; operation = 1'b1; $display("%b", result);

// TEST #221
// -0.0794779755606 - -45.8858072433 = 45.8063292677
// Expected Z = 01000010001101110011100110101110
#10 a = 32'b10111101101000101100010101011001; b = 32'b11000010001101111000101100010001; operation = 1'b1; $display("%b", result);

// TEST #222
// 0.843400829415 - 225.97842275 = -225.13502192
// Expected Z = 11000011011000010010001010010001
#10 a = 32'b00111111010101111110100100011110; b = 32'b01000011011000011111101001111010; operation = 1'b1; $display("%b", result);

// TEST #223
// 0.882835428253 - 203.414682865 = -202.531847436
// Expected Z = 11000011010010101000100000100111
#10 a = 32'b00111111011000100000000110000001; b = 32'b01000011010010110110101000101001; operation = 1'b1; $display("%b", result);

// TEST #224
// -0.0396271122839 + 442.622078725 = 442.582451613
// Expected Z = 01000011110111010100101010001110
#10 a = 32'b10111101001000100101000000001010; b = 32'b01000011110111010100111110100000; operation = 1'b0; $display("%b", result);

// TEST #225
// 0.376164406527 - -276.808837855 = 277.185002261
// Expected Z = 01000011100010101001011110101110
#10 a = 32'b00111110110000001001100010011111; b = 32'b11000011100010100110011110001000; operation = 1'b1; $display("%b", result);

// TEST #226
// 0.67053602057 - -995.804654076 = 996.475190097
// Expected Z = 01000100011110010001111001101010
#10 a = 32'b00111111001010111010100001000000; b = 32'b11000100011110001111001101111111; operation = 1'b1; $display("%b", result);

// TEST #227
// -0.238266470749 + 595.678379498 = 595.440113028
// Expected Z = 01000100000101001101110000101011
#10 a = 32'b10111110011100111111110000100000; b = 32'b01000100000101001110101101101011; operation = 1'b0; $display("%b", result);

// TEST #228
// -0.121265590999 + 805.225915754 = 805.104650163
// Expected Z = 01000100010010010100011010110011
#10 a = 32'b10111101111110000101101000011000; b = 32'b01000100010010010100111001110101; operation = 1'b0; $display("%b", result);

// TEST #229
// 0.383680255122 + 846.532530723 = 846.916210978
// Expected Z = 01000100010100111011101010100011
#10 a = 32'b00111110110001000111000110111101; b = 32'b01000100010100111010001000010101; operation = 1'b0; $display("%b", result);

// TEST #230
// 0.625746285684 - 54.9983966667 = -54.372650381
// Expected Z = 11000010010110010111110110011000
#10 a = 32'b00111111001000000011000011101001; b = 32'b01000010010110111111111001011100; operation = 1'b1; $display("%b", result);

// TEST #231
// 0.300494850145 - 31.6540310502 = -31.3535362001
// Expected Z = 11000001111110101101010000001011
#10 a = 32'b00111110100110011101101001110110; b = 32'b01000001111111010011101101110101; operation = 1'b1; $display("%b", result);

// TEST #232
// -0.791651140139 + 135.890823291 = 135.099172151
// Expected Z = 01000011000001110001100101100011
#10 a = 32'b10111111010010101010100110100110; b = 32'b01000011000001111110010000001101; operation = 1'b0; $display("%b", result);

// TEST #233
// 0.73922334285 - 154.695856669 = -153.956633326
// Expected Z = 11000011000110011111010011100110
#10 a = 32'b00111111001111010011110110111110; b = 32'b01000011000110101011001000100100; operation = 1'b1; $display("%b", result);

// TEST #234
// 0.450258169257 + 637.147064441 = 637.59732261
// Expected Z = 01000100000111110110011000111011
#10 a = 32'b00111110111001101000100000111101; b = 32'b01000100000111110100100101101010; operation = 1'b0; $display("%b", result);

// TEST #235
// -0.536569718023 + -29.4010297137 = -29.9375994317
// Expected Z = 11000001111011111000000000110100
#10 a = 32'b10111111000010010101110010100010; b = 32'b11000001111010110011010101001111; operation = 1'b0; $display("%b", result);

// TEST #236
// -0.155444177778 + -883.488063854 = -883.643508031
// Expected Z = 11000100010111001110100100101111
#10 a = 32'b10111110000111110010110011000010; b = 32'b11000100010111001101111100111100; operation = 1'b0; $display("%b", result);

// TEST #237
// -0.221512644453 + -455.214284148 = -455.435796793
// Expected Z = 11000011111000111011011111001000
#10 a = 32'b10111110011000101101010000110110; b = 32'b11000011111000111001101101101110; operation = 1'b0; $display("%b", result);

// TEST #238
// -0.401798924761 - -122.13436156 = 121.732562635
// Expected Z = 01000010111100110111011100010010
#10 a = 32'b10111110110011011011100010010111; b = 32'b11000010111101000100010011001011; operation = 1'b1; $display("%b", result);

// TEST #239
// -0.683995784689 + 240.03658621 = 239.352590426
// Expected Z = 01000011011011110101101001000011
#10 a = 32'b10111111001011110001101001011001; b = 32'b01000011011100000000100101011110; operation = 1'b0; $display("%b", result);

// TEST #240
// 0.215130112883 - -76.9743851676 = 77.1895152805
// Expected Z = 01000010100110100110000100001000
#10 a = 32'b00111110010111000100101100010001; b = 32'b11000010100110011111001011100011; operation = 1'b1; $display("%b", result);

// TEST #241
// 0.650176137739 + -485.657522133 = -485.007345996
// Expected Z = 11000011111100101000000011110001
#10 a = 32'b00111111001001100111000111110010; b = 32'b11000011111100101101010000101010; operation = 1'b0; $display("%b", result);

// TEST #242
// 0.474122905652 + -99.2413743522 = -98.7672514465
// Expected Z = 11000010110001011000100011010101
#10 a = 32'b00111110111100101100000000111101; b = 32'b11000010110001100111101110010101; operation = 1'b0; $display("%b", result);

// TEST #243
// 0.715967501719 + -981.474883801 = -980.758916299
// Expected Z = 11000100011101010011000010010010
#10 a = 32'b00111111001101110100100110100101; b = 32'b11000100011101010101111001100100; operation = 1'b0; $display("%b", result);

// TEST #244
// -0.143780229458 + -25.0308883695 = -25.174668599
// Expected Z = 11000001110010010110010110111001
#10 a = 32'b10111110000100110011101100100000; b = 32'b11000001110010000011111101000010; operation = 1'b0; $display("%b", result);

// TEST #245
// 0.591383419374 - 470.806570696 = -470.215187277
// Expected Z = 11000011111010110001101110001011
#10 a = 32'b00111111000101110110010011100111; b = 32'b01000011111010110110011100111110; operation = 1'b1; $display("%b", result);

// TEST #246
// -0.817322864036 + 528.213911178 = 527.396588314
// Expected Z = 01000100000000111101100101100010
#10 a = 32'b10111111010100010011110000010010; b = 32'b01000100000001000000110110110001; operation = 1'b0; $display("%b", result);

// TEST #247
// 0.246573589257 + -612.384990494 = -612.138416905
// Expected Z = 11000100000110010000100011011100
#10 a = 32'b00111110011111000111110111001001; b = 32'b11000100000110010001100010100100; operation = 1'b0; $display("%b", result);

// TEST #248
// 0.955226084603 - 801.432544169 = -800.477318085
// Expected Z = 11000100010010000001111010001100
#10 a = 32'b00111111011101001000100110110010; b = 32'b01000100010010000101101110101111; operation = 1'b1; $display("%b", result);

// TEST #249
// 0.580714549493 + 122.466448513 = 123.047163062
// Expected Z = 01000010111101100001100000100110
#10 a = 32'b00111111000101001010100110110101; b = 32'b01000010111101001110111011010010; operation = 1'b0; $display("%b", result);

// TEST #250
// -0.783842289042 - -504.291930736 = 503.508088447
// Expected Z = 01000011111110111100000100001001
#10 a = 32'b10111111010010001010100111100011; b = 32'b11000011111111000010010101011110; operation = 1'b1; $display("%b", result);

// TEST #251
// -0.878708545005 + 112.811814577 = 111.933106032
// Expected Z = 01000010110111111101110111000000
#10 a = 32'b10111111011000001111001100001011; b = 32'b01000010111000011001111110100110; operation = 1'b0; $display("%b", result);

// TEST #252
// -0.550333594937 + 757.730051041 = 757.179717447
// Expected Z = 01000100001111010100101110000000
#10 a = 32'b10111111000011001110001010101010; b = 32'b01000100001111010110111010111001; operation = 1'b0; $display("%b", result);

// TEST #253
// 0.746676769183 + -554.472255957 = -553.725579188
// Expected Z = 11000100000010100110111001110000
#10 a = 32'b00111111001111110010011000110101; b = 32'b11000100000010101001111000111001; operation = 1'b0; $display("%b", result);

// TEST #254
// 0.208232739117 + 555.055240114 = 555.263472853
// Expected Z = 01000100000010101101000011011101
#10 a = 32'b00111110010101010011101011110111; b = 32'b01000100000010101100001110001001; operation = 1'b0; $display("%b", result);

// TEST #255
// 0.746546822528 - -10.8314489426 = 11.5779957651
// Expected Z = 01000001001110010011111101111000
#10 a = 32'b00111111001111110001110110110001; b = 32'b11000001001011010100110110011101; operation = 1'b1; $display("%b", result);

// TEST #256
// -0.575673920982 + 243.662416319 = 243.086742398
// Expected Z = 01000011011100110001011000110101
#10 a = 32'b10111111000100110101111101011110; b = 32'b01000011011100111010100110010100; operation = 1'b0; $display("%b", result);

// TEST #257
// 0.062407674332 + -317.735766751 = -317.673359077
// Expected Z = 11000011100111101101011000110001
#10 a = 32'b00111101011111111001111100110001; b = 32'b11000011100111101101111000101110; operation = 1'b0; $display("%b", result);

// TEST #258
// -0.250755884861 + 261.883741086 = 261.632985201
// Expected Z = 01000011100000101101000100000110
#10 a = 32'b10111110100000000110001100010011; b = 32'b01000011100000101111000100011110; operation = 1'b0; $display("%b", result);

// TEST #259
// -0.0109894341643 - -124.730786191 = 124.719796757
// Expected Z = 01000010111110010111000010001001
#10 a = 32'b10111100001101000000110100000111; b = 32'b11000010111110010111011000101010; operation = 1'b1; $display("%b", result);

// TEST #260
// -0.674369571701 + 200.046290808 = 199.371921237
// Expected Z = 01000011010001110101111100110110
#10 a = 32'b10111111001011001010001101111100; b = 32'b01000011010010000000101111011010; operation = 1'b0; $display("%b", result);

// TEST #261
// 0.716535498189 + -406.936057013 = -406.219521515
// Expected Z = 11000011110010110001110000011001
#10 a = 32'b00111111001101110110111011011111; b = 32'b11000011110010110111011111010001; operation = 1'b0; $display("%b", result);

// TEST #262
// 0.662010828703 + 574.29376785 = 574.955778679
// Expected Z = 01000100000011111011110100101011
#10 a = 32'b00111111001010010111100110001011; b = 32'b01000100000011111001001011001101; operation = 1'b0; $display("%b", result);

// TEST #263
// -0.767313781094 - 654.546637302 = -655.313951083
// Expected Z = 11000100001000111101010000011000
#10 a = 32'b10111111010001000110111010101101; b = 32'b01000100001000111010001011111100; operation = 1'b1; $display("%b", result);

// TEST #264
// 0.692792247516 + 942.014750017 = 942.707542264
// Expected Z = 01000100011010111010110101001000
#10 a = 32'b00111111001100010101101011010101; b = 32'b01000100011010111000000011110010; operation = 1'b0; $display("%b", result);

// TEST #265
// -0.52150926959 - 129.626982448 = -130.148491717
// Expected Z = 11000011000000100010011000000100
#10 a = 32'b10111111000001011000000110100010; b = 32'b01000011000000011010000010000010; operation = 1'b1; $display("%b", result);

// TEST #266
// 0.846251474588 - -822.805473808 = 823.651725282
// Expected Z = 01000100010011011110100110110110
#10 a = 32'b00111111010110001010001111110000; b = 32'b11000100010011011011001110001101; operation = 1'b1; $display("%b", result);

// TEST #267
// 0.382546197091 - -309.896314339 = 310.278860537
// Expected Z = 01000011100110110010001110110010
#10 a = 32'b00111110110000111101110100011000; b = 32'b11000011100110101111001010111010; operation = 1'b1; $display("%b", result);

// TEST #268
// 0.514050115328 - 611.474311282 = -610.960261167
// Expected Z = 11000100000110001011110101110101
#10 a = 32'b00111111000000111001100011001010; b = 32'b01000100000110001101111001011011; operation = 1'b1; $display("%b", result);

// TEST #269
// -0.971112277247 + 813.79501424 = 812.823901962
// Expected Z = 01000100010010110011010010111011
#10 a = 32'b10111111011110001001101011010000; b = 32'b01000100010010110111001011100010; operation = 1'b0; $display("%b", result);

// TEST #270
// 0.684499466263 + 133.967811725 = 134.652311192
// Expected Z = 01000011000001101010011011111110
#10 a = 32'b00111111001011110011101101011011; b = 32'b01000011000001011111011111000011; operation = 1'b0; $display("%b", result);

// TEST #271
// 0.0914988771279 + -168.128064002 = -168.036565125
// Expected Z = 11000011001010000000100101011100
#10 a = 32'b00111101101110110110001111000011; b = 32'b11000011001010000010000011001001; operation = 1'b0; $display("%b", result);

// TEST #272
// 0.0257219853759 + -540.079046358 = -540.053324373
// Expected Z = 11000100000001110000001101101010
#10 a = 32'b00111100110100101011011011101010; b = 32'b11000100000001110000010100001111; operation = 1'b0; $display("%b", result);

// TEST #273
// 0.787020847993 + -904.689249399 = -903.902228551
// Expected Z = 11000100011000011111100110111110
#10 a = 32'b00111111010010010111101000110011; b = 32'b11000100011000100010110000011101; operation = 1'b0; $display("%b", result);

// TEST #274
// 0.29405989182 + 846.022339148 = 846.31639904
// Expected Z = 01000100010100111001010001000000
#10 a = 32'b00111110100101101000111100000101; b = 32'b01000100010100111000000101101110; operation = 1'b0; $display("%b", result);

// TEST #275
// -0.925672796434 - -21.3670704963 = 20.4413976999
// Expected Z = 01000001101000111000011111111100
#10 a = 32'b10111111011011001111100011100100; b = 32'b11000001101010101110111111000011; operation = 1'b1; $display("%b", result);

// TEST #276
// -0.913785269376 - 453.347769319 = -454.261554589
// Expected Z = 11000011111000110010000101111011
#10 a = 32'b10111111011010011110110111010101; b = 32'b01000011111000101010110010000100; operation = 1'b1; $display("%b", result);

// TEST #277
// 0.77586053937 - -149.211043079 = 149.986903618
// Expected Z = 01000011000101011111110010100110
#10 a = 32'b00111111010001101001111011001100; b = 32'b11000011000101010011011000000111; operation = 1'b1; $display("%b", result);

// TEST #278
// 0.885950774305 + -883.440680437 = -882.554729663
// Expected Z = 11000100010111001010001110000001
#10 a = 32'b00111111011000101100110110101100; b = 32'b11000100010111001101110000110100; operation = 1'b0; $display("%b", result);

// TEST #279
// -0.12747428264 + 497.820837525 = 497.693363243
// Expected Z = 01000011111110001101100011000000
#10 a = 32'b10111110000000101000100010011110; b = 32'b01000011111110001110100100010001; operation = 1'b0; $display("%b", result);

// TEST #280
// -0.386545680269 + 416.394201779 = 416.007656098
// Expected Z = 01000011110100000000000011111011
#10 a = 32'b10111110110001011110100101010001; b = 32'b01000011110100000011001001110101; operation = 1'b0; $display("%b", result);

// TEST #281
// 0.864745417721 + 412.832066097 = 413.696811515
// Expected Z = 01000011110011101101100100110001
#10 a = 32'b00111111010111010101111111110101; b = 32'b01000011110011100110101010000001; operation = 1'b0; $display("%b", result);

// TEST #282
// 0.283903147926 - 592.663653059 = -592.379749911
// Expected Z = 11000100000101000001100001001110
#10 a = 32'b00111110100100010101101111000001; b = 32'b01000100000101000010101001111001; operation = 1'b1; $display("%b", result);

// TEST #283
// 0.0040121134374 + 261.357426618 = 261.361438731
// Expected Z = 01000011100000101010111001000100
#10 a = 32'b00111011100000110111100000001100; b = 32'b01000011100000101010110111000000; operation = 1'b0; $display("%b", result);

// TEST #284
// -0.140071069384 + -673.617044145 = -673.757115215
// Expected Z = 11000100001010000111000001110101
#10 a = 32'b10111110000011110110111011001010; b = 32'b11000100001010000110011101111110; operation = 1'b0; $display("%b", result);

// TEST #285
// -0.353131728653 + 231.969461304 = 231.616329575
// Expected Z = 01000011011001111001110111001000
#10 a = 32'b10111110101101001100110110101111; b = 32'b01000011011001111111100000101111; operation = 1'b0; $display("%b", result);

// TEST #286
// -0.991157073252 + -864.517818016 = -865.508975089
// Expected Z = 11000100010110000110000010010011
#10 a = 32'b10111111011111011011110001111000; b = 32'b11000100010110000010000100100100; operation = 1'b0; $display("%b", result);

// TEST #287
// 0.888428362809 + -424.253510574 = -423.365082211
// Expected Z = 11000011110100111010111010111011
#10 a = 32'b00111111011000110111000000001011; b = 32'b11000011110101000010000001110011; operation = 1'b0; $display("%b", result);

// TEST #288
// 0.63447667228 + -379.02022167 = -378.385744998
// Expected Z = 11000011101111010011000101100000
#10 a = 32'b00111111001000100110110100010000; b = 32'b11000011101111011000001010010111; operation = 1'b0; $display("%b", result);

// TEST #289
// 0.718707407592 - 48.5010375029 = -47.7823300953
// Expected Z = 11000010001111110010000100011011
#10 a = 32'b00111111001101111111110100110101; b = 32'b01000010010000100000000100010000; operation = 1'b1; $display("%b", result);

// TEST #290
// 0.94216302166 + -326.923880479 = -325.981717458
// Expected Z = 11000011101000101111110110101001
#10 a = 32'b00111111011100010011000110011001; b = 32'b11000011101000110111011001000010; operation = 1'b0; $display("%b", result);

// TEST #291
// -0.618416334604 + 238.089505483 = 237.471089149
// Expected Z = 01000011011011010111100010011001
#10 a = 32'b10111111000111100101000010001000; b = 32'b01000011011011100001011011101010; operation = 1'b0; $display("%b", result);

// TEST #292
// 0.363530159242 + 340.858336081 = 341.221866241
// Expected Z = 01000011101010101001110001100110
#10 a = 32'b00111110101110100010000010100000; b = 32'b01000011101010100110110111011110; operation = 1'b0; $display("%b", result);

// TEST #293
// 0.18782307625 + -502.860354576 = -502.672531499
// Expected Z = 11000011111110110101011000010110
#10 a = 32'b00111110010000000101010010110001; b = 32'b11000011111110110110111000100000; operation = 1'b0; $display("%b", result);

// TEST #294
// 0.201680245155 + 722.316996351 = 722.518676596
// Expected Z = 01000100001101001010000100110010
#10 a = 32'b00111110010011101000010101000100; b = 32'b01000100001101001001010001001010; operation = 1'b0; $display("%b", result);

// TEST #295
// -0.444068036435 - 863.267953747 = -863.712021783
// Expected Z = 11000100010101111110110110010010
#10 a = 32'b10111110111000110101110011100011; b = 32'b01000100010101111101000100100110; operation = 1'b1; $display("%b", result);

// TEST #296
// 0.646156284633 + 1.08934151149 = 1.73549779612
// Expected Z = 00111111110111100010010011001011
#10 a = 32'b00111111001001010110101010000000; b = 32'b00111111100010110110111110001011; operation = 1'b0; $display("%b", result);

// TEST #297
// -0.1581272726 - 229.946943263 = -230.105070536
// Expected Z = 11000011011001100001101011100110
#10 a = 32'b10111110001000011110110000011110; b = 32'b01000011011001011111001001101011; operation = 1'b1; $display("%b", result);

// TEST #298
// 0.213891501834 - 911.667734051 = -911.45384255
// Expected Z = 11000100011000111101110100001100
#10 a = 32'b00111110010110110000011001100000; b = 32'b01000100011000111110101010111100; operation = 1'b1; $display("%b", result);

// TEST #299
// -0.970973956514 - 962.839139732 = -963.810113689
// Expected Z = 11000100011100001111001111011001
#10 a = 32'b10111111011110001001000111000000; b = 32'b01000100011100001011010110110100; operation = 1'b1; $display("%b", result);

// TEST #300
// -0.696450689907 - -335.945674349 = 335.249223659
// Expected Z = 01000011101001111001111111100111
#10 a = 32'b10111111001100100100101010011000; b = 32'b11000011101001111111100100001100; operation = 1'b1; $display("%b", result);

// TEST #301
// -825253.459132 + -675978.107453 = -1501231.56659
// Expected Z = 11001001101101110100000101111101
#10 a = 32'b11001001010010010111101001010111; b = 32'b11001001001001010000100010100010; operation = 1'b0; $display("%b", result);

// TEST #302
// -519009.093428 + -865712.709781 = -1384721.80321
// Expected Z = 11001001101010010000100010001110
#10 a = 32'b11001000111111010110110000100011; b = 32'b11001001010100110101101100001011; operation = 1'b0; $display("%b", result);

// TEST #303
// -506257.760742 + 486540.912386 = -19716.8483558
// Expected Z = 11000110100110100000100110110010
#10 a = 32'b11001000111101110011001000111000; b = 32'b01001000111011011001000110011101; operation = 1'b0; $display("%b", result);

// TEST #304
// -960380.513116 + -414930.002175 = -1375310.51529
// Expected Z = 11001001101001111110001001110100
#10 a = 32'b11001001011010100111011111001000; b = 32'b11001000110010101001101001000000; operation = 1'b0; $display("%b", result);

// TEST #305
// -928608.196232 - -666677.488359 = -261930.707873
// Expected Z = 11001000011111111100101010101101
#10 a = 32'b11001001011000101011011000000011; b = 32'b11001001001000101100001101011000; operation = 1'b1; $display("%b", result);

// TEST #306
// -191943.933143 - 854228.005311 = -1046171.93845
// Expected Z = 11001001011111110110100110111111
#10 a = 32'b11001000001110110111000111111100; b = 32'b01001001010100001000110101000000; operation = 1'b1; $display("%b", result);

// TEST #307
// 877031.156909 + -845992.005058 = 31039.1518513
// Expected Z = 01000110111100100111111001001110
#10 a = 32'b01001001010101100001111001110011; b = 32'b11001001010011101000101010000000; operation = 1'b0; $display("%b", result);

// TEST #308
// 975673.943168 - -973124.597077 = 1948798.54025
// Expected Z = 01001001111011011110001111110100
#10 a = 32'b01001001011011100011001110011111; b = 32'b11001001011011011001010001001010; operation = 1'b1; $display("%b", result);

// TEST #309
// 619324.006048 - -36871.9715039 = 656195.977552
// Expected Z = 01001001001000000011010001000000
#10 a = 32'b01001001000101110011001111000000; b = 32'b11000111000100000000011111111001; operation = 1'b1; $display("%b", result);

// TEST #310
// -77614.7724777 + -478144.087035 = -555758.859512
// Expected Z = 11001001000001111010111011101110
#10 a = 32'b11000111100101111001011101100011; b = 32'b11001000111010010111100000000011; operation = 1'b0; $display("%b", result);

// TEST #311
// 320213.336929 + -37220.016995 = 282993.319934
// Expected Z = 01001000100010100010111000101010
#10 a = 32'b01001000100111000101101010101011; b = 32'b11000111000100010110010000000100; operation = 1'b0; $display("%b", result);

// TEST #312
// -755909.177105 + 675566.721678 = -80342.4554264
// Expected Z = 11000111100111001110101100111010
#10 a = 32'b11001001001110001000110001010011; b = 32'b01001001001001001110111011101100; operation = 1'b0; $display("%b", result);

// TEST #313
// -518747.115123 - -780439.689632 = 261692.574509
// Expected Z = 01001000011111111000111100100101
#10 a = 32'b11001000111111010100101101100100; b = 32'b11001001001111101000100101111011; operation = 1'b1; $display("%b", result);

// TEST #314
// 519042.660633 - 61900.283293 = 457142.37734
// Expected Z = 01001000110111110011011011001100
#10 a = 32'b01001000111111010111000001010101; b = 32'b01000111011100011100110001001001; operation = 1'b1; $display("%b", result);

// TEST #315
// 107413.545876 - 991829.118514 = -884415.572638
// Expected Z = 11001001010101111110101111111001
#10 a = 32'b01000111110100011100101011000110; b = 32'b01001001011100100010010101010010; operation = 1'b1; $display("%b", result);

// TEST #316
// -548200.521108 + 434451.945819 = -113748.575289
// Expected Z = 11000111110111100010101001001010
#10 a = 32'b11001001000001011101011010001000; b = 32'b01001000110101000010001001111110; operation = 1'b0; $display("%b", result);

// TEST #317
// 898559.634771 + 508814.163794 = 1407373.79856
// Expected Z = 01001001101010111100110001101110
#10 a = 32'b01001001010110110101111111111010; b = 32'b01001000111110000111000111000101; operation = 1'b0; $display("%b", result);

// TEST #318
// 421096.440421 - -147903.478628 = 568999.919049
// Expected Z = 01001001000010101110101001111111
#10 a = 32'b01001000110011011001110100001110; b = 32'b11001000000100000110111111011111; operation = 1'b1; $display("%b", result);

// TEST #319
// -6381.81526538 - -316077.567451 = 309695.752186
// Expected Z = 01001000100101110011011111111000
#10 a = 32'b11000101110001110110111010000110; b = 32'b11001000100110100101010110110010; operation = 1'b1; $display("%b", result);

// TEST #320
// -991976.300078 - 831590.618122 = -1823566.9182
// Expected Z = 11001001110111101001101001110111
#10 a = 32'b11001001011100100010111010000101; b = 32'b01001001010010110000011001101010; operation = 1'b1; $display("%b", result);

// TEST #321
// -412327.783864 - -852872.738894 = 440544.955031
// Expected Z = 01001000110101110001110000011111
#10 a = 32'b11001000110010010101010011111001; b = 32'b11001001010100000011100010001100; operation = 1'b1; $display("%b", result);

// TEST #322
// 475559.096301 + -650203.018619 = -174643.922318
// Expected Z = 11001000001010101000110011111011
#10 a = 32'b01001000111010000011010011100011; b = 32'b11001001000111101011110110110000; operation = 1'b0; $display("%b", result);

// TEST #323
// 106410.211854 - 103935.147489 = 2475.06436505
// Expected Z = 01000101000110101011000100001000
#10 a = 32'b01000111110011111101010100011011; b = 32'b01000111110010101111111110010011; operation = 1'b1; $display("%b", result);

// TEST #324
// 789477.767849 + -842576.885981 = -53099.1181318
// Expected Z = 11000111010011110110101100011110
#10 a = 32'b01001001010000001011111001011100; b = 32'b11001001010011011011010100001110; operation = 1'b0; $display("%b", result);

// TEST #325
// -431956.738057 - -197778.347578 = -234178.390478
// Expected Z = 11001000011001001011000010011001
#10 a = 32'b11001000110100101110101010011000; b = 32'b11001000010000010010010010010110; operation = 1'b1; $display("%b", result);

// TEST #326
// 49961.8732777 + -266804.950397 = -216843.077119
// Expected Z = 11001000010100111100001011000101
#10 a = 32'b01000111010000110010100111100000; b = 32'b11001000100000100100011010011110; operation = 1'b0; $display("%b", result);

// TEST #327
// 513748.536725 - -713684.344592 = 1227432.88132
// Expected Z = 01001001100101011101010101000111
#10 a = 32'b01001000111110101101101010010001; b = 32'b11001001001011100011110101000110; operation = 1'b1; $display("%b", result);

// TEST #328
// -72280.2451371 - 742631.917355 = -814912.162492
// Expected Z = 11001001010001101111010000000011
#10 a = 32'b11000111100011010010110000011111; b = 32'b01001001001101010100111001111111; operation = 1'b1; $display("%b", result);

// TEST #329
// 903933.098462 + 335365.856926 = 1239298.95539
// Expected Z = 01001001100101110100100000011000
#10 a = 32'b01001001010111001010111111010010; b = 32'b01001000101000111100000010111011; operation = 1'b0; $display("%b", result);

// TEST #330
// -584958.102007 - 970530.298565 = -1555488.40057
// Expected Z = 11001001101111011110000100000011
#10 a = 32'b11001001000011101100111111100010; b = 32'b01001001011011001111001000100101; operation = 1'b1; $display("%b", result);

// TEST #331
// 744306.26159 - 280215.396513 = 464090.865076
// Expected Z = 01001000111000101001101101011100
#10 a = 32'b01001001001101011011011100100100; b = 32'b01001000100010001101001011101101; operation = 1'b1; $display("%b", result);

// TEST #332
// -351091.878443 + -16245.0311824 = -367336.909625
// Expected Z = 11001000101100110101110100011101
#10 a = 32'b11001000101010110110111001111100; b = 32'b11000110011111011101010000100000; operation = 1'b0; $display("%b", result);

// TEST #333
// -466499.234372 - 979467.661997 = -1445966.89637
// Expected Z = 11001001101100001000001001110111
#10 a = 32'b11001000111000111100100001100111; b = 32'b01001001011011110010000010111011; operation = 1'b1; $display("%b", result);

// TEST #334
// 255975.661485 - 588308.752899 = -332333.091413
// Expected Z = 11001000101000100100010110100011
#10 a = 32'b01001000011110011111100111101010; b = 32'b01001001000011111010000101001100; operation = 1'b1; $display("%b", result);

// TEST #335
// -587613.487871 + 590573.859122 = 2960.37125083
// Expected Z = 01000101001110010000010111110001
#10 a = 32'b11001001000011110111010111011000; b = 32'b01001001000100000010111011011110; operation = 1'b0; $display("%b", result);

// TEST #336
// 114055.928886 + 320200.622655 = 434256.551541
// Expected Z = 01001000110101000000101000010010
#10 a = 32'b01000111110111101100001111110111; b = 32'b01001000100111000101100100010100; operation = 1'b0; $display("%b", result);

// TEST #337
// 661502.043268 - -178306.285037 = 839808.328306
// Expected Z = 01001001010011010000100000000101
#10 a = 32'b01001001001000010111111111100001; b = 32'b11001000001011100010000010010010; operation = 1'b1; $display("%b", result);

// TEST #338
// 428348.811724 - 557325.984257 = -128977.172533
// Expected Z = 11000111111110111110100010010110
#10 a = 32'b01001000110100010010011110011010; b = 32'b01001001000010000001000011100000; operation = 1'b1; $display("%b", result);

// TEST #339
// 253722.768052 - 92072.2179533 = 161650.550099
// Expected Z = 01001000000111011101110010100011
#10 a = 32'b01001000011101111100011010110001; b = 32'b01000111101100111101010000011100; operation = 1'b1; $display("%b", result);

// TEST #340
// -803938.838497 + -675157.15616 = -1479095.99466
// Expected Z = 11001001101101001000110111000000
#10 a = 32'b11001001010001000100011000101101; b = 32'b11001001001001001101010101010010; operation = 1'b0; $display("%b", result);

// TEST #341
// -334649.106067 - -918540.847559 = 583891.741492
// Expected Z = 01001001000011101000110100111100
#10 a = 32'b11001000101000110110011100100011; b = 32'b11001001011000000100000011001110; operation = 1'b1; $display("%b", result);

// TEST #342
// 56617.4337195 + 235262.752031 = 291880.18575
// Expected Z = 01001000100011101000010100000110
#10 a = 32'b01000111010111010010100101101111; b = 32'b01001000011001011011111110110000; operation = 1'b0; $display("%b", result);

// TEST #343
// -474404.020836 + -670758.112893 = -1145162.13373
// Expected Z = 11001001100010111100101001010001
#10 a = 32'b11001000111001111010010010000001; b = 32'b11001001001000111100001001100010; operation = 1'b0; $display("%b", result);

// TEST #344
// -962813.70477 + 696532.550142 = -266281.154628
// Expected Z = 11001000100000100000010100100101
#10 a = 32'b11001001011010110000111111011011; b = 32'b01001001001010100000110101001001; operation = 1'b0; $display("%b", result);

// TEST #345
// 301311.535773 + 168849.886191 = 470161.421964
// Expected Z = 01001000111001011001001000101110
#10 a = 32'b01001000100100110001111111110001; b = 32'b01001000001001001110010001111001; operation = 1'b0; $display("%b", result);

// TEST #346
// 727404.049032 - -268926.932253 = 996330.981285
// Expected Z = 01001001011100110011111010110000
#10 a = 32'b01001001001100011001011011000001; b = 32'b11001000100000110100111111011110; operation = 1'b1; $display("%b", result);

// TEST #347
// -15531.1277898 + -510805.126066 = -526336.253856
// Expected Z = 11001001000000001000000000000100
#10 a = 32'b11000110011100101010110010000011; b = 32'b11001000111110010110101010100100; operation = 1'b0; $display("%b", result);

// TEST #348
// 222292.365879 - -951266.658678 = 1173559.02456
// Expected Z = 01001001100011110100000110111000
#10 a = 32'b01001000010110010001010100010111; b = 32'b11001001011010000011111000101011; operation = 1'b1; $display("%b", result);

// TEST #349
// -458623.73495 - 946705.375252 = -1405329.1102
// Expected Z = 11001001101010111000110010001001
#10 a = 32'b11001000110111111110111111111000; b = 32'b01001001011001110010000100010110; operation = 1'b1; $display("%b", result);

// TEST #350
// -869425.124572 + 649868.109678 = -219557.014894
// Expected Z = 11001000010101100110100101000001
#10 a = 32'b11001001010101000100001100010010; b = 32'b01001001000111101010100011000010; operation = 1'b0; $display("%b", result);

// TEST #351
// 236714.468102 + 993228.881493 = 1229943.34959
// Expected Z = 01001001100101100010001110111011
#10 a = 32'b01001000011001110010101010011110; b = 32'b01001001011100100111110011001110; operation = 1'b0; $display("%b", result);

// TEST #352
// 935036.836315 + -280531.639155 = 654505.19716
// Expected Z = 01001001000111111100101010010011
#10 a = 32'b01001001011001000100011111001101; b = 32'b11001000100010001111101001110100; operation = 1'b0; $display("%b", result);

// TEST #353
// -277592.301287 - 602625.153684 = -880217.454971
// Expected Z = 11001001010101101110010110010111
#10 a = 32'b11001000100001111000101100001010; b = 32'b01001001000100110010000000010010; operation = 1'b1; $display("%b", result);

// TEST #354
// -251617.947741 + 846477.64941 = 594859.701669
// Expected Z = 01001001000100010011101010111011
#10 a = 32'b11001000011101011011100001111101; b = 32'b01001001010011101010100011011010; operation = 1'b0; $display("%b", result);

// TEST #355
// 326260.932663 - 247505.785744 = 78755.1469199
// Expected Z = 01000111100110011101000110010011
#10 a = 32'b01001000100111110100111010011110; b = 32'b01001000011100011011010001110010; operation = 1'b1; $display("%b", result);

// TEST #356
// -533428.485425 + -94898.8181951 = -628327.30362
// Expected Z = 11001001000110010110011001110101
#10 a = 32'b11001001000000100011101101001000; b = 32'b11000111101110010101100101101001; operation = 1'b0; $display("%b", result);

// TEST #357
// -727986.972831 - 729583.443761 = -1457570.41659
// Expected Z = 11001001101100011110110100010011
#10 a = 32'b11001001001100011011101100110000; b = 32'b01001001001100100001111011110111; operation = 1'b1; $display("%b", result);

// TEST #358
// 562543.857303 - -659014.9245 = 1221558.7818
// Expected Z = 01001001100101010001110110110110
#10 a = 32'b01001001000010010101011011111110; b = 32'b11001001001000001110010001101111; operation = 1'b1; $display("%b", result);

// TEST #359
// -528485.229979 - -515555.693464 = -12929.5365152
// Expected Z = 11000110010010100000011000100101
#10 a = 32'b11001001000000010000011001010100; b = 32'b11001000111110111011110001110110; operation = 1'b1; $display("%b", result);

// TEST #360
// 266333.59694 + 175001.245971 = 441334.842912
// Expected Z = 01001000110101110111111011011011
#10 a = 32'b01001000100000100000101110110011; b = 32'b01001000001010101110011001010000; operation = 1'b0; $display("%b", result);

// TEST #361
// -471135.012553 - 857914.078847 = -1329049.0914
// Expected Z = 11001001101000100011110011001001
#10 a = 32'b11001000111001100000101111100000; b = 32'b01001001010100010111001110100001; operation = 1'b1; $display("%b", result);

// TEST #362
// 130732.726292 + -349092.494543 = -218359.76825
// Expected Z = 11001000010101010011110111110001
#10 a = 32'b01000111111111110101011001011101; b = 32'b11001000101010100111010010010000; operation = 1'b0; $display("%b", result);

// TEST #363
// 267701.177822 - -514069.742782 = 781770.920604
// Expected Z = 01001001001111101101110010101111
#10 a = 32'b01001000100000101011011010100110; b = 32'b11001000111110110000001010111000; operation = 1'b1; $display("%b", result);

// TEST #364
// 6207.21475263 - -328150.694489 = 334357.909241
// Expected Z = 01001000101000110100001010111101
#10 a = 32'b01000101110000011111100110111000; b = 32'b11001000101000000011101011010110; operation = 1'b1; $display("%b", result);

// TEST #365
// 528948.278535 - -561894.81893 = 1090843.09746
// Expected Z = 01001001100001010010100011011001
#10 a = 32'b01001001000000010010001101000100; b = 32'b11001001000010010010111001101101; operation = 1'b1; $display("%b", result);

// TEST #366
// 420404.507138 - 959671.309827 = -539266.802689
// Expected Z = 11001001000000111010100000101101
#10 a = 32'b01001000110011010100011010010000; b = 32'b01001001011010100100101101110101; operation = 1'b1; $display("%b", result);

// TEST #367
// -429619.499056 - 803527.349471 = -1233146.84853
// Expected Z = 11001001100101101000011111010111
#10 a = 32'b11001000110100011100011001110000; b = 32'b01001001010001000010110001110110; operation = 1'b1; $display("%b", result);

// TEST #368
// -761162.021148 - 672505.655507 = -1433667.67666
// Expected Z = 11001001101011110000001000011101
#10 a = 32'b11001001001110011101010010100000; b = 32'b01001001001001000010111110011010; operation = 1'b1; $display("%b", result);

// TEST #369
// 961555.788446 - 772014.074257 = 189541.714189
// Expected Z = 01001000001110010001100101101110
#10 a = 32'b01001001011010101100000100111101; b = 32'b01001001001111000111101011100001; operation = 1'b1; $display("%b", result);

// TEST #370
// 526867.98081 + 912237.635249 = 1439105.61606
// Expected Z = 01001001101011111010110000001101
#10 a = 32'b01001001000000001010000101000000; b = 32'b01001001010111101011011011011010; operation = 1'b0; $display("%b", result);

// TEST #371
// -43895.8452896 - -814301.883631 = 770406.038341
// Expected Z = 01001001001111000001011001100001
#10 a = 32'b11000111001010110111011111011000; b = 32'b11001001010001101100110111011110; operation = 1'b1; $display("%b", result);

// TEST #372
// 839680.456584 + 531999.249283 = 1371679.70587
// Expected Z = 01001001101001110111000011111110
#10 a = 32'b01001001010011010000000000000111; b = 32'b01001001000000011110000111110100; operation = 1'b0; $display("%b", result);

// TEST #373
// 84666.6547997 - 753165.59566 = -668498.940861
// Expected Z = 11001001001000110011010100101111
#10 a = 32'b01000111101001010101110101010100; b = 32'b01001001001101111110000011011010; operation = 1'b1; $display("%b", result);

// TEST #374
// 234257.101349 + -642867.070975 = -408609.969626
// Expected Z = 11001000110001111000010000111111
#10 a = 32'b01001000011001001100010001000110; b = 32'b11001001000111001111001100110001; operation = 1'b0; $display("%b", result);

// TEST #375
// -114112.315093 + -973759.092445 = -1087871.40754
// Expected Z = 11001001100001001100101111111011
#10 a = 32'b11000111110111101110000000101000; b = 32'b11001001011011011011101111110001; operation = 1'b0; $display("%b", result);

// TEST #376
// 290067.41069 + 237574.722963 = 527642.133653
// Expected Z = 01001001000000001101000110100010
#10 a = 32'b01001000100011011010001001101101; b = 32'b01001000011010000000000110101110; operation = 1'b0; $display("%b", result);

// TEST #377
// -760841.992307 - 22229.0889453 = -783071.081252
// Expected Z = 11001001001111110010110111110001
#10 a = 32'b11001001001110011100000010100000; b = 32'b01000110101011011010101000101110; operation = 1'b1; $display("%b", result);

// TEST #378
// -21697.7353455 - 350806.951256 = -372504.686601
// Expected Z = 11001000101101011110001100010110
#10 a = 32'b11000110101010011000001101111000; b = 32'b01001000101010110100101011011110; operation = 1'b1; $display("%b", result);

// TEST #379
// 51860.5359832 - 923027.431453 = -871166.89547
// Expected Z = 11001001010101001010111111101110
#10 a = 32'b01000111010010101001010010001001; b = 32'b01001001011000010101100100110111; operation = 1'b1; $display("%b", result);

// TEST #380
// 694250.516094 - 944245.257071 = -249994.740977
// Expected Z = 11001000011101000010001010101111
#10 a = 32'b01001001001010010111111010101000; b = 32'b01001001011001101000011101010100; operation = 1'b1; $display("%b", result);

// TEST #381
// 165250.325608 + 231292.496612 = 396542.82222
// Expected Z = 01001000110000011001111111011010
#10 a = 32'b01001000001000010110000010010101; b = 32'b01001000011000011101111100100000; operation = 1'b0; $display("%b", result);

// TEST #382
// -800697.855743 - -193999.709566 = -606698.146177
// Expected Z = 11001001000101000001111010100010
#10 a = 32'b11001001010000110111101110011110; b = 32'b11001000001111010111001111101101; operation = 1'b1; $display("%b", result);

// TEST #383
// 897725.640765 + 668620.913809 = 1566346.55457
// Expected Z = 01001001101111110011010001010100
#10 a = 32'b01001001010110110010101111011010; b = 32'b01001001001000110011110011001111; operation = 1'b0; $display("%b", result);

// TEST #384
// 880915.162757 + 28590.8822469 = 909506.045004
// Expected Z = 01001001010111100000110000100001
#10 a = 32'b01001001010101110001000100110011; b = 32'b01000110110111110101110111000100; operation = 1'b0; $display("%b", result);

// TEST #385
// 105568.317119 - -288686.051933 = 394254.369052
// Expected Z = 01001000110000001000000111001100
#10 a = 32'b01000111110011100011000000101001; b = 32'b11001000100011001111010111000010; operation = 1'b1; $display("%b", result);

// TEST #386
// 678956.803978 + -630267.391854 = 48689.412124
// Expected Z = 01000111001111100011000101101010
#10 a = 32'b01001001001001011100001011001101; b = 32'b11001001000110011101111110110110; operation = 1'b0; $display("%b", result);

// TEST #387
// -334311.610387 + -496737.818379 = -831049.428766
// Expected Z = 11001001010010101110010010010111
#10 a = 32'b11001000101000110011110011110100; b = 32'b11001000111100101000110000111010; operation = 1'b0; $display("%b", result);

// TEST #388
// -747917.062199 + -798695.792721 = -1546612.85492
// Expected Z = 11001001101111001100101110100111
#10 a = 32'b11001001001101101001100011010001; b = 32'b11001001010000101111111001111101; operation = 1'b0; $display("%b", result);

// TEST #389
// -326701.37176 + 312660.251047 = -14041.1207137
// Expected Z = 11000110010110110110010001111100
#10 a = 32'b11001000100111111000010110101100; b = 32'b01001000100110001010101010001000; operation = 1'b0; $display("%b", result);

// TEST #390
// 541221.827664 - -961276.556008 = 1502498.38367
// Expected Z = 01001001101101110110100100010011
#10 a = 32'b01001001000001000010001001011101; b = 32'b11001001011010101010111111001001; operation = 1'b1; $display("%b", result);

// TEST #391
// 245879.565407 + 377625.745523 = 623505.31093
// Expected Z = 01001001000110000011100100010101
#10 a = 32'b01001000011100000001110111100100; b = 32'b01001000101110000110001100111000; operation = 1'b0; $display("%b", result);

// TEST #392
// 16363.5727819 + -391761.094552 = -375397.52177
// Expected Z = 11001000101101110100110010110001
#10 a = 32'b01000110011111111010111001001011; b = 32'b11001000101111110100101000100011; operation = 1'b0; $display("%b", result);

// TEST #393
// -56525.3382007 + 780169.477812 = 723644.139611
// Expected Z = 01001001001100001010101111000010
#10 a = 32'b11000111010111001100110101010111; b = 32'b01001001001111100111100010011000; operation = 1'b0; $display("%b", result);

// TEST #394
// 602782.43246 + 135633.839517 = 738416.271978
// Expected Z = 01001001001101000100011100000100
#10 a = 32'b01001001000100110010100111100111; b = 32'b01001000000001000111010001110110; operation = 1'b0; $display("%b", result);

// TEST #395
// 329253.076463 - 323668.664726 = 5584.41173742
// Expected Z = 01000101101011101000001101001011
#10 a = 32'b01001000101000001100010010100010; b = 32'b01001000100111100000101010010101; operation = 1'b1; $display("%b", result);

// TEST #396
// -941510.894466 + 71429.8002831 = -870081.094183
// Expected Z = 11001001010101000110110000010010
#10 a = 32'b11001001011001011101110001101110; b = 32'b01000111100010111000001011100110; operation = 1'b0; $display("%b", result);

// TEST #397
// 523683.448862 + 442569.259215 = 966252.708077
// Expected Z = 01001001011010111110011011001011
#10 a = 32'b01001000111111111011010001101110; b = 32'b01001000110110000001100100101000; operation = 1'b0; $display("%b", result);

// TEST #398
// 45396.1591053 + -117579.974691 = -72183.8155857
// Expected Z = 11000111100011001111101111101000
#10 a = 32'b01000111001100010101010000101001; b = 32'b11000111111001011010010111111101; operation = 1'b0; $display("%b", result);

// TEST #399
// -941333.936813 - -93733.3954931 = -847600.54132
// Expected Z = 11001001010011101110111100001001
#10 a = 32'b11001001011001011101000101011111; b = 32'b11000111101101110001001010110011; operation = 1'b1; $display("%b", result);

// TEST #400
// -205211.346557 + 21324.6465411 = -183886.700016
// Expected Z = 11001000001100111001001110101101
#10 a = 32'b11001000010010000110011011010110; b = 32'b01000110101001101001100101001011; operation = 1'b0; $display("%b", result);

// TEST #401
// 215.561299749 + -0.796808026434 = 214.764491723
// Expected Z = 01000011010101101100001110110110
#10 a = 32'b01000011010101111000111110110001; b = 32'b10111111010010111111101110011100; operation = 1'b0; $display("%b", result);

// TEST #402
// -741.333801914 + 0.725506396311 = -740.608295518
// Expected Z = 11000100001110010010011011101110
#10 a = 32'b11000100001110010101010101011101; b = 32'b00111111001110011011101011001010; operation = 1'b0; $display("%b", result);

// TEST #403
// 313.334496504 + -0.584240903023 = 312.750255601
// Expected Z = 01000011100111000110000000001000
#10 a = 32'b01000011100111001010101011010001; b = 32'b10111111000101011001000011010000; operation = 1'b0; $display("%b", result);

// TEST #404
// -138.18455512 + -0.988249190606 = -139.172804311
// Expected Z = 11000011000010110010110000111101
#10 a = 32'b11000011000010100010111100111111; b = 32'b10111111011111001111110111100110; operation = 1'b0; $display("%b", result);

// TEST #405
// -387.143829036 - 0.129077952083 = -387.272906988
// Expected Z = 11000011110000011010001011101111
#10 a = 32'b11000011110000011001001001101001; b = 32'b00111110000001000010110100000011; operation = 1'b1; $display("%b", result);

// TEST #406
// -377.378587433 - 0.244893910083 = -377.623481343
// Expected Z = 11000011101111001100111111001110
#10 a = 32'b11000011101111001011000001110110; b = 32'b00111110011110101100010101111000; operation = 1'b1; $display("%b", result);

// TEST #407
// -539.748292541 - 0.80386388533 = -540.552156426
// Expected Z = 11000100000001110010001101010111
#10 a = 32'b11000100000001101110111111100100; b = 32'b00111111010011011100101000000110; operation = 1'b1; $display("%b", result);

// TEST #408
// 776.044209737 - -0.894398241285 = 776.938607978
// Expected Z = 01000100010000100011110000010010
#10 a = 32'b01000100010000100000001011010100; b = 32'b10111111011001001111011101001000; operation = 1'b1; $display("%b", result);

// TEST #409
// -217.804904688 + -0.860052743912 = -218.664957431
// Expected Z = 11000011010110101010101000111011
#10 a = 32'b11000011010110011100111000001110; b = 32'b10111111010111000010110001101011; operation = 1'b0; $display("%b", result);

// TEST #410
// 88.0951131001 + -0.421187553176 = 87.673925547
// Expected Z = 01000010101011110101100100001101
#10 a = 32'b01000010101100000011000010110011; b = 32'b10111110110101111010010111100101; operation = 1'b0; $display("%b", result);

// TEST #411
// 724.421339295 + -0.0499470909951 = 724.371392204
// Expected Z = 01000100001101010001011111000101
#10 a = 32'b01000100001101010001101011110111; b = 32'b10111101010011001001010101010010; operation = 1'b0; $display("%b", result);

// TEST #412
// -581.124326855 + -0.687308410851 = -581.811635266
// Expected Z = 11000100000100010111001111110010
#10 a = 32'b11000100000100010100011111110101; b = 32'b10111111001011111111001101110010; operation = 1'b0; $display("%b", result);

// TEST #413
// -197.535898117 - 0.737798723311 = -198.27369684
// Expected Z = 11000011010001100100011000010001
#10 a = 32'b11000011010001011000100100110001; b = 32'b00111111001111001110000001100001; operation = 1'b1; $display("%b", result);

// TEST #414
// 144.398278155 - 0.920430832995 = 143.477847322
// Expected Z = 01000011000011110111101001010100
#10 a = 32'b01000011000100000110010111110110; b = 32'b00111111011010111010000101011011; operation = 1'b1; $display("%b", result);

// TEST #415
// 16.9687833065 - 0.382374727299 = 16.5864085792
// Expected Z = 01000001100001001011000011110111
#10 a = 32'b01000001100001111100000000010001; b = 32'b00111110110000111100011010011111; operation = 1'b1; $display("%b", result);

// TEST #416
// 535.999488952 - -0.15638478899 = 536.155873741
// Expected Z = 01000100000001100000100111111010
#10 a = 32'b01000100000001011111111111111000; b = 32'b10111110001000000010001101010110; operation = 1'b1; $display("%b", result);

// TEST #417
// 911.655391766 - -0.73203099028 = 912.387422756
// Expected Z = 01000100011001000001100011001100
#10 a = 32'b01000100011000111110100111110010; b = 32'b10111111001110110110011001100010; operation = 1'b1; $display("%b", result);

// TEST #418
// -193.181614795 - 0.488637541387 = -193.670252336
// Expected Z = 11000011010000011010101110010110
#10 a = 32'b11000011010000010010111001111110; b = 32'b00111110111110100010111010110011; operation = 1'b1; $display("%b", result);

// TEST #419
// 877.815554418 - 0.492433220289 = 877.323121198
// Expected Z = 01000100010110110101010010101110
#10 a = 32'b01000100010110110111010000110010; b = 32'b00111110111111000010000000110101; operation = 1'b1; $display("%b", result);

// TEST #420
// 352.182584905 + -0.268331036716 = 351.914253869
// Expected Z = 01000011101011111111010100000110
#10 a = 32'b01000011101100000001011101011111; b = 32'b10111110100010010110001010110000; operation = 1'b0; $display("%b", result);

// TEST #421
// -849.222314158 + -0.966856255668 = -850.189170413
// Expected Z = 11000100010101001000110000011011
#10 a = 32'b11000100010101000100111000111010; b = 32'b10111111011101111000001111100100; operation = 1'b0; $display("%b", result);

// TEST #422
// -310.514743545 + 0.918779664221 = -309.595963881
// Expected Z = 11000011100110101100110001001001
#10 a = 32'b11000011100110110100000111100011; b = 32'b00111111011010110011010100100101; operation = 1'b0; $display("%b", result);

// TEST #423
// -87.8579574874 - -0.0425989365155 = -87.8153585508
// Expected Z = 11000010101011111010000101110111
#10 a = 32'b11000010101011111011011101000110; b = 32'b10111101001011100111110000111001; operation = 1'b1; $display("%b", result);

// TEST #424
// 93.7440134974 - 0.772068701445 = 92.971944796
// Expected Z = 01000010101110011111000110100011
#10 a = 32'b01000010101110110111110011101111; b = 32'b00111111010001011010011001001011; operation = 1'b1; $display("%b", result);

// TEST #425
// 121.140575561 + -0.632411484602 = 120.508164077
// Expected Z = 01000010111100010000010000101110
#10 a = 32'b01000010111100100100011111111010; b = 32'b10111111001000011110010110111000; operation = 1'b0; $display("%b", result);

// TEST #426
// 962.773372331 - -0.667506289311 = 963.44087862
// Expected Z = 01000100011100001101110000110111
#10 a = 32'b01000100011100001011000101111111; b = 32'b10111111001010101110000110110001; operation = 1'b1; $display("%b", result);

// TEST #427
// -851.354478143 + 0.874335373274 = -850.48014277
// Expected Z = 11000100010101001001111010111011
#10 a = 32'b11000100010101001101011010110000; b = 32'b00111111010111111101010001110001; operation = 1'b0; $display("%b", result);

// TEST #428
// 726.594172874 - 0.60582087932 = 725.988351995
// Expected Z = 01000100001101010111111101000001
#10 a = 32'b01000100001101011010011000000111; b = 32'b00111111000110110001011100010100; operation = 1'b1; $display("%b", result);

// TEST #429
// -320.219621245 + -0.730291459803 = -320.949912705
// Expected Z = 11000011101000000111100110010111
#10 a = 32'b11000011101000000001110000011101; b = 32'b10111111001110101111010001100010; operation = 1'b0; $display("%b", result);

// TEST #430
// -607.400599983 + -0.00802951532639 = -607.408629498
// Expected Z = 11000100000101111101101000100111
#10 a = 32'b11000100000101111101100110100011; b = 32'b10111100000000111000111000111010; operation = 1'b0; $display("%b", result);

// TEST #431
// -125.65674741 - 0.758809696281 = -126.415557107
// Expected Z = 11000010111111001101010011000100
#10 a = 32'b11000010111110110101000001000001; b = 32'b00111111010000100100000101011010; operation = 1'b1; $display("%b", result);

// TEST #432
// 478.769564607 - -0.832909030347 = 479.602473638
// Expected Z = 01000011111011111100110100011110
#10 a = 32'b01000011111011110110001010000001; b = 32'b10111111010101010011100110000111; operation = 1'b1; $display("%b", result);

// TEST #433
// 463.68415792 + -0.479505481484 = 463.204652439
// Expected Z = 01000011111001111001101000110010
#10 a = 32'b01000011111001111101011110010010; b = 32'b10111110111101011000000110111110; operation = 1'b0; $display("%b", result);

// TEST #434
// -496.101592734 + 0.206563303149 = -495.895029431
// Expected Z = 11000011111101111111001010010000
#10 a = 32'b11000011111110000000110100000001; b = 32'b00111110010100111000010101010101; operation = 1'b0; $display("%b", result);

// TEST #435
// 484.750789202 - -0.506636411734 = 485.257425614
// Expected Z = 01000011111100101010000011110011
#10 a = 32'b01000011111100100110000000011010; b = 32'b10111111000000011011001011101101; operation = 1'b1; $display("%b", result);

// TEST #436
// 342.418738477 + 0.171219231694 = 342.589957709
// Expected Z = 01000011101010110100101110000100
#10 a = 32'b01000011101010110011010110011001; b = 32'b00111110001011110101010000011000; operation = 1'b0; $display("%b", result);

// TEST #437
// -19.5756345415 + -0.715376605016 = -20.2910111465
// Expected Z = 11000001101000100101001111111110
#10 a = 32'b11000001100111001001101011100110; b = 32'b10111111001101110010001011101100; operation = 1'b0; $display("%b", result);

// TEST #438
// 601.214733951 - -0.148287890249 = 601.363021841
// Expected Z = 01000100000101100101011100111100
#10 a = 32'b01000100000101100100110110111110; b = 32'b10111110000101111101100011001000; operation = 1'b1; $display("%b", result);

// TEST #439
// -572.478927236 + -0.697184406094 = -573.176111642
// Expected Z = 11000100000011110100101101000101
#10 a = 32'b11000100000011110001111010100111; b = 32'b10111111001100100111101010101101; operation = 1'b0; $display("%b", result);

// TEST #440
// 487.610320196 + 0.114004055192 = 487.724324251
// Expected Z = 01000011111100111101110010110111
#10 a = 32'b01000011111100111100111000011111; b = 32'b00111101111010010111101011110101; operation = 1'b0; $display("%b", result);

// TEST #441
// -853.959593921 + 0.706310230393 = -853.253283691
// Expected Z = 11000100010101010101000000110110
#10 a = 32'b11000100010101010111110101101010; b = 32'b00111111001101001101000010111111; operation = 1'b0; $display("%b", result);

// TEST #442
// 522.117670384 - -0.981445314637 = 523.099115699
// Expected Z = 01000100000000101100011001011000
#10 a = 32'b01000100000000101000011110001000; b = 32'b10111111011110110100000000000000; operation = 1'b1; $display("%b", result);

// TEST #443
// -765.738924418 - 0.244739336474 = -765.983663755
// Expected Z = 11000100001111110111111011110100
#10 a = 32'b11000100001111110110111101001011; b = 32'b00111110011110101001110011110011; operation = 1'b1; $display("%b", result);

// TEST #444
// 161.626138915 + -0.173833369306 = 161.452305546
// Expected Z = 01000011001000010111001111001010
#10 a = 32'b01000011001000011010000001001011; b = 32'b10111110001100100000000101100000; operation = 1'b0; $display("%b", result);

// TEST #445
// -571.894161887 + 0.0136986325894 = -571.880463255
// Expected Z = 11000100000011101111100001011010
#10 a = 32'b11000100000011101111100100111010; b = 32'b00111100011000000111000000111011; operation = 1'b0; $display("%b", result);

// TEST #446
// 870.859088118 - -0.106136426009 = 870.965224544
// Expected Z = 01000100010110011011110111000110
#10 a = 32'b01000100010110011011011011111011; b = 32'b10111101110110010101111000001110; operation = 1'b1; $display("%b", result);

// TEST #447
// 309.360288209 - 0.855282063201 = 308.505006146
// Expected Z = 01000011100110100100000010100100
#10 a = 32'b01000011100110101010111000011110; b = 32'b00111111010110101111001111000100; operation = 1'b1; $display("%b", result);

// TEST #448
// -699.643848085 + -0.383011184068 = -700.026859269
// Expected Z = 11000100001011110000000110111000
#10 a = 32'b11000100001011101110100100110101; b = 32'b10111110110001000001101000001011; operation = 1'b0; $display("%b", result);

// TEST #449
// -146.56725907 + -0.936889169184 = -147.50414824
// Expected Z = 11000011000100111000000100010000
#10 a = 32'b11000011000100101001000100111000; b = 32'b10111111011011111101011111111000; operation = 1'b0; $display("%b", result);

// TEST #450
// -217.316043526 + 0.791773226726 = -216.524270299
// Expected Z = 11000011010110001000011000110111
#10 a = 32'b11000011010110010101000011101000; b = 32'b00111111010010101011000110100110; operation = 1'b0; $display("%b", result);

// TEST #451
// 396.752825348 + 0.54021059879 = 397.293035947
// Expected Z = 01000011110001101010010110000010
#10 a = 32'b01000011110001100110000001011101; b = 32'b00111111000010100100101100111110; operation = 1'b0; $display("%b", result);

// TEST #452
// -957.535647423 + -0.182646662744 = -957.718294086
// Expected Z = 11000100011011110110110111111001
#10 a = 32'b11000100011011110110001001001000; b = 32'b10111110001110110000011110111010; operation = 1'b0; $display("%b", result);

// TEST #453
// -106.015278779 - -0.243834785163 = -105.771443994
// Expected Z = 11000010110100111000101011111011
#10 a = 32'b11000010110101000000011111010011; b = 32'b10111110011110011010111111010011; operation = 1'b1; $display("%b", result);

// TEST #454
// 78.1624522202 + 0.169081844897 = 78.3315340651
// Expected Z = 01000010100111001010100110111111
#10 a = 32'b01000010100111000101001100101101; b = 32'b00111110001011010010001111001011; operation = 1'b0; $display("%b", result);

// TEST #455
// -69.9201045082 + -0.971373991622 = -70.8914784998
// Expected Z = 11000010100011011100100001110000
#10 a = 32'b11000010100010111101011100011000; b = 32'b10111111011110001010101111110111; operation = 1'b0; $display("%b", result);

// TEST #456
// 463.098709861 - 0.427452213558 = 462.671257648
// Expected Z = 01000011111001110101010111101100
#10 a = 32'b01000011111001111000110010100011; b = 32'b00111110110110101101101100000100; operation = 1'b1; $display("%b", result);

// TEST #457
// -824.943814582 - 0.927948374152 = -825.871762956
// Expected Z = 11000100010011100111011111001011
#10 a = 32'b11000100010011100011110001100111; b = 32'b00111111011011011000111000000110; operation = 1'b1; $display("%b", result);

// TEST #458
// 986.499802903 - 0.0369319427886 = 986.46287096
// Expected Z = 01000100011101101001110110100000
#10 a = 32'b01000100011101101001111111111101; b = 32'b00111101000101110100010111110011; operation = 1'b1; $display("%b", result);

// TEST #459
// 769.813983072 - -0.78688866903 = 770.600871741
// Expected Z = 01000100010000001010011001110101
#10 a = 32'b01000100010000000111010000011000; b = 32'b10111111010010010111000110001001; operation = 1'b1; $display("%b", result);

// TEST #460
// 8.40543105421 - 0.820148529799 = 7.58528252441
// Expected Z = 01000000111100101011101010100010
#10 a = 32'b01000001000001100111110010100101; b = 32'b00111111010100011111010101000001; operation = 1'b1; $display("%b", result);

// TEST #461
// -391.751034584 + 0.890069633574 = -390.860964951
// Expected Z = 11000011110000110110111000110100
#10 a = 32'b11000011110000111110000000100010; b = 32'b00111111011000111101101110011010; operation = 1'b0; $display("%b", result);

// TEST #462
// -69.141105274 + 0.884693494928 = -68.2564117791
// Expected Z = 11000010100010001000001101001000
#10 a = 32'b11000010100010100100100000111111; b = 32'b00111111011000100111101101000110; operation = 1'b0; $display("%b", result);

// TEST #463
// 804.973045901 + -0.872698441548 = 804.100347459
// Expected Z = 01000100010010010000011001101100
#10 a = 32'b01000100010010010011111001000110; b = 32'b10111111010111110110100100101010; operation = 1'b0; $display("%b", result);

// TEST #464
// -193.595289221 + -0.517914017323 = -194.113203239
// Expected Z = 11000011010000100001110011111011
#10 a = 32'b11000011010000011001100001100101; b = 32'b10111111000001001001011000000011; operation = 1'b0; $display("%b", result);

// TEST #465
// -930.002874052 + -0.968611901997 = -930.971485954
// Expected Z = 11000100011010001011111000101101
#10 a = 32'b11000100011010001000000000101111; b = 32'b10111111011101111111011011110011; operation = 1'b0; $display("%b", result);

// TEST #466
// 740.983647978 + 0.36369980742 = 741.347347785
// Expected Z = 01000100001110010101011000111011
#10 a = 32'b01000100001110010011111011110100; b = 32'b00111110101110100011011011011100; operation = 1'b0; $display("%b", result);

// TEST #467
// -523.680556819 - -0.0781767596907 = -523.602380059
// Expected Z = 11000100000000101110011010001101
#10 a = 32'b11000100000000101110101110001110; b = 32'b10111101101000000001101100100011; operation = 1'b1; $display("%b", result);

// TEST #468
// -355.375068378 + 0.463788423371 = -354.911279955
// Expected Z = 11000011101100010111010010100101
#10 a = 32'b11000011101100011011000000000010; b = 32'b00111110111011010111010110101101; operation = 1'b0; $display("%b", result);

// TEST #469
// -403.48640296 + -0.0949548716839 = -403.581357831
// Expected Z = 11000011110010011100101001101010
#10 a = 32'b11000011110010011011111001000010; b = 32'b10111101110000100111011110110011; operation = 1'b0; $display("%b", result);

// TEST #470
// -897.958409186 + -0.174696774422 = -898.13310596
// Expected Z = 11000100011000001000100010000101
#10 a = 32'b11000100011000000111110101010111; b = 32'b10111110001100101110001110110110; operation = 1'b0; $display("%b", result);

// TEST #471
// -145.763989299 - 0.339471706813 = -146.103461005
// Expected Z = 11000011000100100001101001111100
#10 a = 32'b11000011000100011100001110010101; b = 32'b00111110101011011100111100111100; operation = 1'b1; $display("%b", result);

// TEST #472
// -701.14809528 - 0.265846859579 = -701.41394214
// Expected Z = 11000100001011110101101001111110
#10 a = 32'b11000100001011110100100101111010; b = 32'b00111110100010000001110100010100; operation = 1'b1; $display("%b", result);

// TEST #473
// 844.845263303 - 0.800070413113 = 844.045192889
// Expected Z = 01000100010100110000001011100100
#10 a = 32'b01000100010100110011011000011001; b = 32'b00111111010011001101000101101010; operation = 1'b1; $display("%b", result);

// TEST #474
// 569.128167187 - -0.643287073132 = 569.77145426
// Expected Z = 01000100000011100111000101100000
#10 a = 32'b01000100000011100100100000110100; b = 32'b10111111001001001010111001110110; operation = 1'b1; $display("%b", result);

// TEST #475
// -673.205548526 - 0.718736574806 = -673.924285101
// Expected Z = 11000100001010000111101100100111
#10 a = 32'b11000100001010000100110100101000; b = 32'b00111111001101111111111100011111; operation = 1'b1; $display("%b", result);

// TEST #476
// -430.197956523 + 0.727985404382 = -429.469971119
// Expected Z = 11000011110101101011110000101000
#10 a = 32'b11000011110101110001100101010111; b = 32'b00111111001110100101110101000000; operation = 1'b0; $display("%b", result);

// TEST #477
// 405.185194517 + 0.203621728126 = 405.388816245
// Expected Z = 01000011110010101011000111000101
#10 a = 32'b01000011110010101001011110110100; b = 32'b00111110010100001000001000110111; operation = 1'b0; $display("%b", result);

// TEST #478
// -611.614621974 - -0.332311568552 = -611.282310405
// Expected Z = 11000100000110001101001000010001
#10 a = 32'b11000100000110001110011101010110; b = 32'b10111110101010100010010010111110; operation = 1'b1; $display("%b", result);

// TEST #479
// 316.471779085 + 0.608724123797 = 317.080503209
// Expected Z = 01000011100111101000101001001110
#10 a = 32'b01000011100111100011110001100011; b = 32'b00111111000110111101010101011000; operation = 1'b0; $display("%b", result);

// TEST #480
// 832.140583169 + -0.838005282814 = 831.302577886
// Expected Z = 01000100010011111101001101011101
#10 a = 32'b01000100010100000000100011111111; b = 32'b10111111010101101000011110000100; operation = 1'b0; $display("%b", result);

// TEST #481
// -272.40857956 - -0.882322060933 = -271.526257499
// Expected Z = 11000011100001111100001101011100
#10 a = 32'b11000011100010000011010001001100; b = 32'b10111111011000011101111111011100; operation = 1'b1; $display("%b", result);

// TEST #482
// -936.695148389 + 0.996483397113 = -935.698664992
// Expected Z = 11000100011010011110110010110111
#10 a = 32'b11000100011010100010110001111101; b = 32'b00111111011111110001100110001001; operation = 1'b0; $display("%b", result);

// TEST #483
// -941.800356088 + -0.500946300727 = -942.301302388
// Expected Z = 11000100011010111001001101001001
#10 a = 32'b11000100011010110111001100111001; b = 32'b10111111000000000011111000000100; operation = 1'b0; $display("%b", result);

// TEST #484
// -793.940582696 + 0.32223007946 = -793.618352617
// Expected Z = 11000100010001100110011110010011
#10 a = 32'b11000100010001100111110000110011; b = 32'b00111110101001001111101101010111; operation = 1'b0; $display("%b", result);

// TEST #485
// 620.820062736 - 0.576546466151 = 620.24351627
// Expected Z = 01000100000110110000111110010110
#10 a = 32'b01000100000110110011010001111100; b = 32'b00111111000100111001100010001101; operation = 1'b1; $display("%b", result);

// TEST #486
// -182.77233245 - -0.609944633616 = -182.162387817
// Expected Z = 11000011001101100010100110010010
#10 a = 32'b11000011001101101100010110111000; b = 32'b10111111000111000010010101010101; operation = 1'b1; $display("%b", result);

// TEST #487
// 938.378535055 + 0.0659746950892 = 938.44450975
// Expected Z = 01000100011010101001110001110011
#10 a = 32'b01000100011010101001100000111010; b = 32'b00111101100001110001110110111110; operation = 1'b0; $display("%b", result);

// TEST #488
// -542.741203537 + -0.723533570223 = -543.464737107
// Expected Z = 11000100000001111101110110111110
#10 a = 32'b11000100000001111010111101110000; b = 32'b10111111001110010011100101111111; operation = 1'b0; $display("%b", result);

// TEST #489
// -692.190404249 + -0.966534796118 = -693.156939045
// Expected Z = 11000100001011010100101000001011
#10 a = 32'b11000100001011010000110000110000; b = 32'b10111111011101110110111011010011; operation = 1'b0; $display("%b", result);

// TEST #490
// -141.157659032 - -0.226178720588 = -140.931480312
// Expected Z = 11000011000011001110111001110101
#10 a = 32'b11000011000011010010100001011100; b = 32'b10111110011001111001101101100101; operation = 1'b1; $display("%b", result);

// TEST #491
// -848.523948106 + -0.0264342611398 = -848.550382367
// Expected Z = 11000100010101000010001100111001
#10 a = 32'b11000100010101000010000110001000; b = 32'b10111100110110001000110010101010; operation = 1'b0; $display("%b", result);

// TEST #492
// -410.791446888 - 0.295707550993 = -411.087154439
// Expected Z = 11000011110011011000101100101000
#10 a = 32'b11000011110011010110010101001110; b = 32'b00111110100101110110011011111011; operation = 1'b1; $display("%b", result);

// TEST #493
// -118.175501832 + 0.466212967046 = -117.709288865
// Expected Z = 11000010111010110110101100101000
#10 a = 32'b11000010111011000101100111011011; b = 32'b00111110111011101011001101110111; operation = 1'b0; $display("%b", result);

// TEST #494
// 902.078889556 + 0.468714259501 = 902.547603816
// Expected Z = 01000100011000011010001100001100
#10 a = 32'b01000100011000011000010100001101; b = 32'b00111110111011111111101101010001; operation = 1'b0; $display("%b", result);

// TEST #495
// 809.520881194 + 0.64962915516 = 810.170510349
// Expected Z = 01000100010010101000101011101010
#10 a = 32'b01000100010010100110000101010110; b = 32'b00111111001001100100111000011001; operation = 1'b0; $display("%b", result);

// TEST #496
// 222.790737397 - -0.379116237536 = 223.169853634
// Expected Z = 01000011010111110010101101111100
#10 a = 32'b01000011010111101100101001101110; b = 32'b10111110110000100001101110000110; operation = 1'b1; $display("%b", result);

// TEST #497
// -507.424829547 + -0.153604358134 = -507.578433905
// Expected Z = 11000011111111011100101000001010
#10 a = 32'b11000011111111011011011001100001; b = 32'b10111110000111010100101001110110; operation = 1'b0; $display("%b", result);

// TEST #498
// 196.794164678 + 0.943223805056 = 197.737388483
// Expected Z = 01000011010001011011110011000101
#10 a = 32'b01000011010001001100101101001110; b = 32'b00111111011100010111011100011110; operation = 1'b0; $display("%b", result);

// TEST #499
// -276.363768589 + 0.303176711277 = -276.060591877
// Expected Z = 11000011100010100000011111000001
#10 a = 32'b11000011100010100010111010010000; b = 32'b00111110100110110011100111111010; operation = 1'b0; $display("%b", result);

// TEST #500
// 30.615877866 + 0.436840924949 = 31.0527187909
// Expected Z = 01000001111110000110101111111000
#10 a = 32'b01000001111101001110110101010001; b = 32'b00111110110111111010100110011101; operation = 1'b0; $display("%b", result);

// TEST #501
// -380040.351591 - -0.0399990036279 = -380040.311592
// Expected Z = 11001000101110011001000100001010
#10 a = 32'b11001000101110011001000100001011; b = 32'b10111101001000111101010111111111; operation = 1'b1; $display("%b", result);

// TEST #502
// -877809.594729 - 0.0244713310668 = -877809.6192
// Expected Z = 11001001010101100100111100011010
#10 a = 32'b11001001010101100100111100011010; b = 32'b00111100110010000111100000011010; operation = 1'b1; $display("%b", result);

// TEST #503
// -160257.457375 - 0.0660339773438 = -160257.523409
// Expected Z = 11001000000111001000000001100001
#10 a = 32'b11001000000111001000000001011101; b = 32'b00111101100001110011110011010010; operation = 1'b1; $display("%b", result);

// TEST #504
// -270688.510356 + -0.0413607060311 = -270688.551717
// Expected Z = 11001000100001000010110000010010
#10 a = 32'b11001000100001000010110000010000; b = 32'b10111101001010010110100111011000; operation = 1'b0; $display("%b", result);

// TEST #505
// -244568.644414 - 0.0716636750627 = -244568.716078
// Expected Z = 11001000011011101101011000101110
#10 a = 32'b11001000011011101101011000101001; b = 32'b00111101100100101100010001101000; operation = 1'b1; $display("%b", result);

// TEST #506
// 150426.86881 + -0.0457079657237 = 150426.823102
// Expected Z = 01001000000100101110011010110101
#10 a = 32'b01001000000100101110011010111000; b = 32'b10111101001110110011100001000111; operation = 1'b0; $display("%b", result);

// TEST #507
// 909254.982566 + 0.00786408278188 = 909254.99043
// Expected Z = 01001001010111011111110001110000
#10 a = 32'b01001001010111011111110001110000; b = 32'b00111100000000001101100001011011; operation = 1'b0; $display("%b", result);

// TEST #508
// 840200.563955 + 0.0100838118235 = 840200.574039
// Expected Z = 01001001010011010010000010001001
#10 a = 32'b01001001010011010010000010001001; b = 32'b00111100001001010011011010010011; operation = 1'b0; $display("%b", result);

// TEST #509
// -324128.116313 - -0.0826026782596 = -324128.033711
// Expected Z = 11001000100111100100010000000001
#10 a = 32'b11001000100111100100010000000100; b = 32'b10111101101010010010101110011000; operation = 1'b1; $display("%b", result);

// TEST #510
// -16076.3506724 - 0.0779185359762 = -16076.4285909
// Expected Z = 11000110011110110011000110110111
#10 a = 32'b11000110011110110011000101100111; b = 32'b00111101100111111001001111000001; operation = 1'b1; $display("%b", result);

// TEST #511
// -86121.6510392 + 0.090585047757 = -86121.5604542
// Expected Z = 11000111101010000011010011001000
#10 a = 32'b11000111101010000011010011010011; b = 32'b00111101101110011000010010100111; operation = 1'b0; $display("%b", result);

// TEST #512
// -33841.0249864 - -0.0550422463597 = -33840.9699442
// Expected Z = 11000111000001000011000011111000
#10 a = 32'b11000111000001000011000100000110; b = 32'b10111101011000010111001111111011; operation = 1'b1; $display("%b", result);

// TEST #513
// -389609.135743 + 0.0688798899612 = -389609.066863
// Expected Z = 11001000101111100011110100100010
#10 a = 32'b11001000101111100011110100100100; b = 32'b00111101100011010001000011100110; operation = 1'b0; $display("%b", result);

// TEST #514
// 335786.004619 + -0.0781229361117 = 335785.926496
// Expected Z = 01001000101000111111010100111110
#10 a = 32'b01001000101000111111010101000000; b = 32'b10111101100111111111111011101011; operation = 1'b0; $display("%b", result);

// TEST #515
// 958173.141465 - -0.0833766222357 = 958173.224842
// Expected Z = 01001001011010011110110111010100
#10 a = 32'b01001001011010011110110111010010; b = 32'b10111101101010101100000101011101; operation = 1'b1; $display("%b", result);

// TEST #516
// 626040.081166 - -0.0322456478957 = 626040.113412
// Expected Z = 01001001000110001101011110000010
#10 a = 32'b01001001000110001101011110000001; b = 32'b10111101000001000001010000000011; operation = 1'b1; $display("%b", result);

// TEST #517
// -585880.857305 + -0.043833561708 = -585880.901139
// Expected Z = 11001001000011110000100110001110
#10 a = 32'b11001001000011110000100110001110; b = 32'b10111101001100111000101011010010; operation = 1'b0; $display("%b", result);

// TEST #518
// 593917.735881 + -0.0109841042634 = 593917.724897
// Expected Z = 01001001000100001111111111011100
#10 a = 32'b01001001000100001111111111011100; b = 32'b10111100001100111111011010101100; operation = 1'b0; $display("%b", result);

// TEST #519
// -420396.453797 + -0.0367955713289 = -420396.490593
// Expected Z = 11001000110011010100010110010000
#10 a = 32'b11001000110011010100010110001111; b = 32'b10111101000101101011011011110100; operation = 1'b0; $display("%b", result);

// TEST #520
// 164766.014125 - -0.0333905236086 = 164766.047515
// Expected Z = 01001000001000001110011110000011
#10 a = 32'b01001000001000001110011110000001; b = 32'b10111101000010001100010010000000; operation = 1'b1; $display("%b", result);

// TEST #521
// -543846.930958 + 0.045958062607 = -543846.885
// Expected Z = 11001001000001001100011001101110
#10 a = 32'b11001001000001001100011001101111; b = 32'b00111101001111000011111010000101; operation = 1'b0; $display("%b", result);

// TEST #522
// 616996.46137 - 0.0389277637179 = 616996.422442
// Expected Z = 01001001000101101010001001000111
#10 a = 32'b01001001000101101010001001000111; b = 32'b00111101000111110111001010111000; operation = 1'b1; $display("%b", result);

// TEST #523
// 522054.096886 - -0.0678903989638 = 522054.164777
// Expected Z = 01001000111111101110100011000101
#10 a = 32'b01001000111111101110100011000011; b = 32'b10111101100010110000101000011111; operation = 1'b1; $display("%b", result);

// TEST #524
// 468669.346677 + -0.0124517572715 = 468669.334225
// Expected Z = 01001000111001001101011110101011
#10 a = 32'b01001000111001001101011110101011; b = 32'b10111100010011000000001001110101; operation = 1'b0; $display("%b", result);

// TEST #525
// 313457.785106 + -0.0539799766185 = 313457.731126
// Expected Z = 01001000100110010000111000110111
#10 a = 32'b01001000100110010000111000111001; b = 32'b10111101010111010001101000011100; operation = 1'b0; $display("%b", result);

// TEST #526
// 104698.551784 + -0.0811308967344 = 104698.470653
// Expected Z = 01000111110011000111110100111100
#10 a = 32'b01000111110011000111110101000111; b = 32'b10111101101001100010011111110101; operation = 1'b0; $display("%b", result);

// TEST #527
// -51517.7441075 + -0.0381779666438 = -51517.7822855
// Expected Z = 11000111010010010011110111001000
#10 a = 32'b11000111010010010011110110111110; b = 32'b10111101000111000110000010000000; operation = 1'b0; $display("%b", result);

// TEST #528
// 864458.9919 + 0.0383061104622 = 864459.030206
// Expected Z = 01001001010100110000110010110000
#10 a = 32'b01001001010100110000110010110000; b = 32'b00111101000111001110011011011110; operation = 1'b0; $display("%b", result);

// TEST #529
// 262485.889564 + 0.00809891508161 = 262485.897663
// Expected Z = 01001000100000000010101010111101
#10 a = 32'b01001000100000000010101010111100; b = 32'b00111100000001001011000101010000; operation = 1'b0; $display("%b", result);

// TEST #530
// 167012.330146 + -0.0415223432576 = 167012.288624
// Expected Z = 01001000001000110001100100010010
#10 a = 32'b01001000001000110001100100010101; b = 32'b10111101001010100001001101010101; operation = 1'b0; $display("%b", result);

// TEST #531
// -425520.989713 + 0.0988988688449 = -425520.890814
// Expected Z = 11001000110011111100011000011101
#10 a = 32'b11001000110011111100011000100000; b = 32'b00111101110010101000101101111101; operation = 1'b0; $display("%b", result);

// TEST #532
// 848796.183207 - 0.0277538452571 = 848796.155453
// Expected Z = 01001001010011110011100111000010
#10 a = 32'b01001001010011110011100111000011; b = 32'b00111100111000110101110000001000; operation = 1'b1; $display("%b", result);

// TEST #533
// 364836.992503 + 0.0553534292992 = 364837.047857
// Expected Z = 01001000101100100010010010100010
#10 a = 32'b01001000101100100010010010100000; b = 32'b00111101011000101011101001000111; operation = 1'b0; $display("%b", result);

// TEST #534
// 257432.490293 + 0.0495198263333 = 257432.539813
// Expected Z = 01001000011110110110011000100011
#10 a = 32'b01001000011110110110011000011111; b = 32'b00111101010010101101010101001101; operation = 1'b0; $display("%b", result);

// TEST #535
// 75451.9082784 - -0.0920109666576 = 75452.0002894
// Expected Z = 01000111100100110101111000000000
#10 a = 32'b01000111100100110101110111110100; b = 32'b10111101101111000111000000111111; operation = 1'b1; $display("%b", result);

// TEST #536
// 544676.104807 + 0.0757523533254 = 544676.180559
// Expected Z = 01001001000001001111101001000011
#10 a = 32'b01001001000001001111101001000010; b = 32'b00111101100110110010010000001101; operation = 1'b0; $display("%b", result);

// TEST #537
// -136185.838894 - 0.0185070403842 = -136185.857401
// Expected Z = 11001000000001001111111001110111
#10 a = 32'b11001000000001001111111001110110; b = 32'b00111100100101111001110000010100; operation = 1'b1; $display("%b", result);

// TEST #538
// -257615.582762 - -0.0977169891595 = -257615.485045
// Expected Z = 11001000011110111001001111011111
#10 a = 32'b11001000011110111001001111100101; b = 32'b10111101110010000001111111011000; operation = 1'b1; $display("%b", result);

// TEST #539
// 699373.445133 - 0.0299139471439 = 699373.415219
// Expected Z = 01001001001010101011111011010111
#10 a = 32'b01001001001010101011111011010111; b = 32'b00111100111101010000111000011000; operation = 1'b1; $display("%b", result);

// TEST #540
// -110798.619979 + -0.071289848347 = -110798.691269
// Expected Z = 11000111110110000110011101011000
#10 a = 32'b11000111110110000110011101001111; b = 32'b10111101100100100000000001101001; operation = 1'b0; $display("%b", result);

// TEST #541
// -183025.365581 + 0.0788608955621 = -183025.28672
// Expected Z = 11001000001100101011110001010010
#10 a = 32'b11001000001100101011110001010111; b = 32'b00111101101000011000000111010010; operation = 1'b0; $display("%b", result);

// TEST #542
// -160548.024488 - -0.0465077743194 = -160547.977981
// Expected Z = 11001000000111001100100011111111
#10 a = 32'b11001000000111001100100100000010; b = 32'b10111101001111100111111011110000; operation = 1'b1; $display("%b", result);

// TEST #543
// 475021.978367 - -0.0383826904851 = 475022.01675
// Expected Z = 01001000111001111111000111000001
#10 a = 32'b01001000111001111111000110111111; b = 32'b10111101000111010011011100101011; operation = 1'b1; $display("%b", result);

// TEST #544
// -85097.538893 - -0.00659240608178 = -85097.5323006
// Expected Z = 11000111101001100011010011000100
#10 a = 32'b11000111101001100011010011000101; b = 32'b10111011110110000000010100011100; operation = 1'b1; $display("%b", result);

// TEST #545
// -214755.373496 - 0.00467140544453 = -214755.378167
// Expected Z = 11001000010100011011100011011000
#10 a = 32'b11001000010100011011100011011000; b = 32'b00111011100110010001001010010111; operation = 1'b1; $display("%b", result);

// TEST #546
// -973782.824452 - 0.0996708346973 = -973782.924123
// Expected Z = 11001001011011011011110101101111
#10 a = 32'b11001001011011011011110101101101; b = 32'b00111101110011000010000000111001; operation = 1'b1; $display("%b", result);

// TEST #547
// -763255.043075 - 0.0760715161024 = -763255.119146
// Expected Z = 11001001001110100101011101110010
#10 a = 32'b11001001001110100101011101110001; b = 32'b00111101100110111100101101100010; operation = 1'b1; $display("%b", result);

// TEST #548
// 935410.738721 - -0.0475137878481 = 935410.786235
// Expected Z = 01001001011001000101111100101101
#10 a = 32'b01001001011001000101111100101100; b = 32'b10111101010000101001110111010001; operation = 1'b1; $display("%b", result);

// TEST #549
// 637354.213529 + -0.0343990427074 = 637354.17913
// Expected Z = 01001001000110111001101010100011
#10 a = 32'b01001001000110111001101010100011; b = 32'b10111101000011001110011000000011; operation = 1'b0; $display("%b", result);

// TEST #550
// -455869.579231 + -0.0855985642884 = -455869.66483
// Expected Z = 11001000110111101001011110110101
#10 a = 32'b11001000110111101001011110110011; b = 32'b10111101101011110100111001001101; operation = 1'b0; $display("%b", result);

// TEST #551
// -350247.686414 - 0.0615287010184 = -350247.747943
// Expected Z = 11001000101010110000010011111000
#10 a = 32'b11001000101010110000010011110110; b = 32'b00111101011111000000010110000101; operation = 1'b1; $display("%b", result);

// TEST #552
// -866536.755391 - -0.00845319048507 = -866536.746938
// Expected Z = 11001001010100111000111010001100
#10 a = 32'b11001001010100111000111010001100; b = 32'b10111100000010100111111101000000; operation = 1'b1; $display("%b", result);

// TEST #553
// -768088.733146 + -0.0954658008358 = -768088.828612
// Expected Z = 11001001001110111000010110001101
#10 a = 32'b11001001001110111000010110001100; b = 32'b10111101110000111000001110010011; operation = 1'b0; $display("%b", result);

// TEST #554
// -69578.3080847 + -0.0650687696827 = -69578.3731535
// Expected Z = 11000111100001111110010100110000
#10 a = 32'b11000111100001111110010100100111; b = 32'b10111101100001010100001011000110; operation = 1'b0; $display("%b", result);

// TEST #555
// -916044.982809 - 0.00213874165251 = -916044.984947
// Expected Z = 11001001010111111010010011010000
#10 a = 32'b11001001010111111010010011010000; b = 32'b00111011000011000010101000100001; operation = 1'b1; $display("%b", result);

// TEST #556
// -320174.179618 + 0.0325216892878 = -320174.147096
// Expected Z = 11001000100111000101010111000101
#10 a = 32'b11001000100111000101010111000110; b = 32'b00111101000001010011010101110110; operation = 1'b0; $display("%b", result);

// TEST #557
// -239481.132979 - 0.0480266008266 = -239481.181006
// Expected Z = 11001000011010011101111001001100
#10 a = 32'b11001000011010011101111001001001; b = 32'b00111101010001001011011110001010; operation = 1'b1; $display("%b", result);

// TEST #558
// -885432.410907 - -0.0690827236556 = -885432.341824
// Expected Z = 11001001010110000010101110000101
#10 a = 32'b11001001010110000010101110000111; b = 32'b10111101100011010111101100111110; operation = 1'b1; $display("%b", result);

// TEST #559
// 482576.03823 - 0.0854443976823 = 482575.952786
// Expected Z = 01001000111010111010000111111110
#10 a = 32'b01001000111010111010001000000001; b = 32'b00111101101011101111110101111001; operation = 1'b1; $display("%b", result);

// TEST #560
// -583323.027503 + -0.0291564667203 = -583323.056659
// Expected Z = 11001001000011100110100110110001
#10 a = 32'b11001001000011100110100110110000; b = 32'b10111100111011101101100110001011; operation = 1'b0; $display("%b", result);

// TEST #561
// 303685.721129 - 0.0844932220595 = 303685.636636
// Expected Z = 01001000100101000100100010110100
#10 a = 32'b01001000100101000100100010110111; b = 32'b00111101101011010000101011001000; operation = 1'b1; $display("%b", result);

// TEST #562
// 725742.135636 - 0.0352425664578 = 725742.100394
// Expected Z = 01001001001100010010111011100010
#10 a = 32'b01001001001100010010111011100010; b = 32'b00111101000100000101101010000010; operation = 1'b1; $display("%b", result);

// TEST #563
// -342022.684606 + 0.059388878501 = -342022.625217
// Expected Z = 11001000101001110000000011010100
#10 a = 32'b11001000101001110000000011010110; b = 32'b00111101011100110100000111000001; operation = 1'b0; $display("%b", result);

// TEST #564
// 84655.9119654 - 0.00841146999022 = 84655.903554
// Expected Z = 01000111101001010101011111110100
#10 a = 32'b01000111101001010101011111110101; b = 32'b00111100000010011101000001000011; operation = 1'b1; $display("%b", result);

// TEST #565
// 856303.906397 - -0.0805557633097 = 856303.986953
// Expected Z = 01001001010100010000111100000000
#10 a = 32'b01001001010100010000111011111111; b = 32'b10111101101001001111101001101100; operation = 1'b1; $display("%b", result);

// TEST #566
// 765814.799363 - 0.0481200890423 = 765814.751243
// Expected Z = 01001001001110101111011101101100
#10 a = 32'b01001001001110101111011101101101; b = 32'b00111101010001010001100110010010; operation = 1'b1; $display("%b", result);

// TEST #567
// 326951.891545 - -0.0476048594855 = 326951.939149
// Expected Z = 01001000100111111010010011111110
#10 a = 32'b01001000100111111010010011111101; b = 32'b10111101010000101111110101010000; operation = 1'b1; $display("%b", result);

// TEST #568
// 864492.130048 - 0.023108559297 = 864492.10694
// Expected Z = 01001001010100110000111011000010
#10 a = 32'b01001001010100110000111011000010; b = 32'b00111100101111010100111000101001; operation = 1'b1; $display("%b", result);

// TEST #569
// 366027.999719 + -0.0498369512888 = 366027.949882
// Expected Z = 01001000101100101011100101111110
#10 a = 32'b01001000101100101011100110000000; b = 32'b10111101010011000010000111010101; operation = 1'b0; $display("%b", result);

// TEST #570
// -529421.26454 + 0.0155132308752 = -529421.249026
// Expected Z = 11001001000000010100000011010100
#10 a = 32'b11001001000000010100000011010100; b = 32'b00111100011111100010101100110101; operation = 1'b0; $display("%b", result);

// TEST #571
// 764200.516739 - 0.0548755970207 = 764200.461864
// Expected Z = 01001001001110101001001010000111
#10 a = 32'b01001001001110101001001010001000; b = 32'b00111101011000001100010100111100; operation = 1'b1; $display("%b", result);

// TEST #572
// 41342.2525227 - -0.0175009801235 = 41342.2700236
// Expected Z = 01000111001000010111111001000101
#10 a = 32'b01000111001000010111111001000001; b = 32'b10111100100011110101111000110111; operation = 1'b1; $display("%b", result);

// TEST #573
// -556884.072021 + 0.0464119270299 = -556884.025609
// Expected Z = 11001001000001111111010101000000
#10 a = 32'b11001001000001111111010101000001; b = 32'b00111101001111100001101001101111; operation = 1'b0; $display("%b", result);

// TEST #574
// 394363.42445 - -0.0425106088103 = 394363.46696
// Expected Z = 01001000110000001000111101101111
#10 a = 32'b01001000110000001000111101101110; b = 32'b10111101001011100001111110011011; operation = 1'b1; $display("%b", result);

// TEST #575
// 70070.4809362 - 0.00611191346016 = 70070.4748243
// Expected Z = 01000111100010001101101100111101
#10 a = 32'b01000111100010001101101100111110; b = 32'b00111011110010000100011001110010; operation = 1'b1; $display("%b", result);

// TEST #576
// -55352.0607505 - -0.00552744747021 = -55352.0552231
// Expected Z = 11000111010110000011100000001110
#10 a = 32'b11000111010110000011100000010000; b = 32'b10111011101101010001111110010111; operation = 1'b1; $display("%b", result);

// TEST #577
// 206080.475273 - 0.0003481743393 = 206080.474924
// Expected Z = 01001000010010010100000000011110
#10 a = 32'b01001000010010010100000000011110; b = 32'b00111001101101101000101100101011; operation = 1'b1; $display("%b", result);

// TEST #578
// 643311.759392 + 0.0978079733784 = 643311.8572
// Expected Z = 01001001000111010000111011111110
#10 a = 32'b01001001000111010000111011111100; b = 32'b00111101110010000100111110001100; operation = 1'b0; $display("%b", result);

// TEST #579
// 192460.961797 - -0.0742805036969 = 192461.036077
// Expected Z = 01001000001110111111001101000010
#10 a = 32'b01001000001110111111001100111110; b = 32'b10111101100110000010000001100000; operation = 1'b1; $display("%b", result);

// TEST #580
// -891367.844645 + 0.0295111720297 = -891367.815134
// Expected Z = 11001001010110011001111001111101
#10 a = 32'b11001001010110011001111001111110; b = 32'b00111100111100011100000101101010; operation = 1'b0; $display("%b", result);

// TEST #581
// 32849.2730571 + -0.0256487683751 = 32849.2474084
// Expected Z = 01000111000000000101000100111111
#10 a = 32'b01000111000000000101000101000110; b = 32'b10111100110100100001110101011110; operation = 1'b0; $display("%b", result);

// TEST #582
// -878975.816533 - 0.00819847568838 = -878975.824732
// Expected Z = 11001001010101101001011111111101
#10 a = 32'b11001001010101101001011111111101; b = 32'b00111100000001100101001011100110; operation = 1'b1; $display("%b", result);

// TEST #583
// 731280.577151 + -0.0227281503566 = 731280.554422
// Expected Z = 01001001001100101000100100001001
#10 a = 32'b01001001001100101000100100001001; b = 32'b10111100101110100011000001100011; operation = 1'b0; $display("%b", result);

// TEST #584
// -708349.871138 + -0.081332161593 = -708349.95247
// Expected Z = 11001001001011001110111111011111
#10 a = 32'b11001001001011001110111111011110; b = 32'b10111101101001101001000101111010; operation = 1'b0; $display("%b", result);

// TEST #585
// 287932.791884 - -0.0722405243441 = 287932.864124
// Expected Z = 01001000100011001001011110011100
#10 a = 32'b01001000100011001001011110011001; b = 32'b10111101100100111111001011010111; operation = 1'b1; $display("%b", result);

// TEST #586
// 474468.993202 + -0.0171863699239 = 474468.976016
// Expected Z = 01001000111001111010110010011111
#10 a = 32'b01001000111001111010110010100000; b = 32'b10111100100011001100101001101110; operation = 1'b0; $display("%b", result);

// TEST #587
// 266087.974821 + 0.00949812845825 = 266087.98432
// Expected Z = 01001000100000011110110011111111
#10 a = 32'b01001000100000011110110011111111; b = 32'b00111100000110111001111000001010; operation = 1'b0; $display("%b", result);

// TEST #588
// -647274.346544 + -0.0224972945081 = -647274.369041
// Expected Z = 11001001000111100000011010100110
#10 a = 32'b11001001000111100000011010100110; b = 32'b10111100101110000100110000111111; operation = 1'b0; $display("%b", result);

// TEST #589
// 996136.161188 - 0.0192582167793 = 996136.14193
// Expected Z = 01001001011100110011001010000010
#10 a = 32'b01001001011100110011001010000011; b = 32'b00111100100111011100001101101000; operation = 1'b1; $display("%b", result);

// TEST #590
// -542239.648573 + -0.0146201451453 = -542239.663193
// Expected Z = 11001001000001000110000111111011
#10 a = 32'b11001001000001000110000111111010; b = 32'b10111100011011111000100101010101; operation = 1'b0; $display("%b", result);

// TEST #591
// 117434.721277 - -0.00803111831113 = 117434.729309
// Expected Z = 01000111111001010101110101011101
#10 a = 32'b01000111111001010101110101011100; b = 32'b10111100000000111001010011110100; operation = 1'b1; $display("%b", result);

// TEST #592
// -29903.7606061 - 0.0687453681465 = -29903.8293514
// Expected Z = 11000110111010011001111110101001
#10 a = 32'b11000110111010011001111110000101; b = 32'b00111101100011001100101001011111; operation = 1'b1; $display("%b", result);

// TEST #593
// 449803.145206 - 0.0859347126082 = 449803.059271
// Expected Z = 01001000110110111010000101100010
#10 a = 32'b01001000110110111010000101100101; b = 32'b00111101101011111111111010001010; operation = 1'b1; $display("%b", result);

// TEST #594
// 855150.502929 + 0.0959665303094 = 855150.598895
// Expected Z = 01001001010100001100011011101010
#10 a = 32'b01001001010100001100011011101000; b = 32'b00111101110001001000101000011010; operation = 1'b0; $display("%b", result);

// TEST #595
// -42952.1015961 - -0.0715322551433 = -42952.0300638
// Expected Z = 11000111001001111100100000001000
#10 a = 32'b11000111001001111100100000011010; b = 32'b10111101100100100111111110000001; operation = 1'b1; $display("%b", result);

// TEST #596
// -451944.95167 - -0.0999228343 = -451944.851748
// Expected Z = 11001000110111001010110100011011
#10 a = 32'b11001000110111001010110100011110; b = 32'b10111101110011001010010001011000; operation = 1'b1; $display("%b", result);

// TEST #597
// -990251.879558 + 0.010403370184 = -990251.869155
// Expected Z = 11001001011100011100001010111110
#10 a = 32'b11001001011100011100001010111110; b = 32'b00111100001010100111001011100110; operation = 1'b0; $display("%b", result);

// TEST #598
// 392690.18375 + 0.0544271921213 = 392690.238177
// Expected Z = 01001000101111111011111001001000
#10 a = 32'b01001000101111111011111001000110; b = 32'b00111101010111101110111100001100; operation = 1'b0; $display("%b", result);

// TEST #599
// -586050.114973 + 0.0799299587893 = -586050.035043
// Expected Z = 11001001000011110001010000100001
#10 a = 32'b11001001000011110001010000100010; b = 32'b00111101101000111011001001010001; operation = 1'b0; $display("%b", result);

// TEST #600
// -486508.997705 - -0.0290665535647 = -486508.968638
// Expected Z = 11001000111011011000110110011111
#10 a = 32'b11001000111011011000110110100000; b = 32'b10111100111011100001110011111011; operation = 1'b1; $display("%b", result);

// TEST #601
// 488247.140211 + 2.00466840938e-06 = 488247.140213
// Expected Z = 01001000111011100110011011100100
#10 a = 32'b01001000111011100110011011100100; b = 32'b00110110000001101000011111110001; operation = 1'b0; $display("%b", result);

// TEST #602
// -391491.553407 - -0.000706155264592 = -391491.552701
// Expected Z = 11001000101111110010100001110010
#10 a = 32'b11001000101111110010100001110010; b = 32'b10111010001110010001110101000111; operation = 1'b1; $display("%b", result);

// TEST #603
// 122425.525038 - 8.29619953045e-07 = 122425.525037
// Expected Z = 01000111111011110001110011000011
#10 a = 32'b01000111111011110001110011000011; b = 32'b00110101010111101011001100001101; operation = 1'b1; $display("%b", result);

// TEST #604
// 355449.69737 + 0.000369887449787 = 355449.69774
// Expected Z = 01001000101011011000111100110110
#10 a = 32'b01001000101011011000111100110110; b = 32'b00111001110000011110110101110100; operation = 1'b0; $display("%b", result);

// TEST #605
// -444316.104683 + 0.000458512027044 = -444316.104225
// Expected Z = 11001000110110001111001110000011
#10 a = 32'b11001000110110001111001110000011; b = 32'b00111001111100000110010001110001; operation = 1'b0; $display("%b", result);

// TEST #606
// 285527.101638 + 0.000345833892633 = 285527.101984
// Expected Z = 01001000100010110110101011100011
#10 a = 32'b01001000100010110110101011100011; b = 32'b00111001101101010101000100001010; operation = 1'b0; $display("%b", result);

// TEST #607
// -120234.865749 + 0.000620471648187 = -120234.865129
// Expected Z = 11000111111010101101010101101111
#10 a = 32'b11000111111010101101010101101111; b = 32'b00111010001000101010011100100110; operation = 1'b0; $display("%b", result);

// TEST #608
// 161999.787904 + 0.000387788402525 = 161999.788292
// Expected Z = 01001000000111100011001111110010
#10 a = 32'b01001000000111100011001111110010; b = 32'b00111001110010110101000000010100; operation = 1'b0; $display("%b", result);

// TEST #609
// 982652.847772 - 8.66325119241e-05 = 982652.847685
// Expected Z = 01001001011011111110011111001110
#10 a = 32'b01001001011011111110011111001110; b = 32'b00111000101101011010111001111010; operation = 1'b1; $display("%b", result);

// TEST #610
// 477000.68837 - 1.76419886776e-05 = 477000.688352
// Expected Z = 01001000111010001110100100010110
#10 a = 32'b01001000111010001110100100010110; b = 32'b00110111100100111111110111100010; operation = 1'b1; $display("%b", result);

// TEST #611
// 696229.010579 + 0.000701015482108 = 696229.01128
// Expected Z = 01001001001010011111101001010000
#10 a = 32'b01001001001010011111101001010000; b = 32'b00111010001101111100010001011010; operation = 1'b0; $display("%b", result);

// TEST #612
// -216849.694152 + -0.000328325229391 = -216849.69448
// Expected Z = 11001000010100111100010001101100
#10 a = 32'b11001000010100111100010001101100; b = 32'b10111001101011000010001100010001; operation = 1'b0; $display("%b", result);

// TEST #613
// -256780.00692 - -0.000738349488197 = -256780.006182
// Expected Z = 11001000011110101100001100000000
#10 a = 32'b11001000011110101100001100000000; b = 32'b10111010010000011000110111001100; operation = 1'b1; $display("%b", result);

// TEST #614
// 452617.493392 - -0.000544206179112 = 452617.493936
// Expected Z = 01001000110111010000000100110000
#10 a = 32'b01001000110111010000000100110000; b = 32'b10111010000011101010100100001111; operation = 1'b1; $display("%b", result);

// TEST #615
// 889157.577973 - -0.000946433345411 = 889157.57892
// Expected Z = 01001001010110010001010001011001
#10 a = 32'b01001001010110010001010001011001; b = 32'b10111010011110000001101000010001; operation = 1'b1; $display("%b", result);

// TEST #616
// 155693.06651 + -0.000885037416541 = 155693.065625
// Expected Z = 01001000000110000000101101000100
#10 a = 32'b01001000000110000000101101000100; b = 32'b10111010011010000000000111011011; operation = 1'b0; $display("%b", result);

// TEST #617
// 144699.511476 + -0.000302096420416 = 144699.511174
// Expected Z = 01001000000011010100111011100001
#10 a = 32'b01001000000011010100111011100001; b = 32'b10111001100111100110001010110010; operation = 1'b0; $display("%b", result);

// TEST #618
// 39780.5818203 + -0.000276050197476 = 39780.5815442
// Expected Z = 01000111000110110110010010010101
#10 a = 32'b01000111000110110110010010010101; b = 32'b10111001100100001011101011010101; operation = 1'b0; $display("%b", result);

// TEST #619
// -477424.308088 - -0.000367832943014 = -477424.30772
// Expected Z = 11001000111010010001111000001010
#10 a = 32'b11001000111010010001111000001010; b = 32'b10111001110000001101100110110100; operation = 1'b1; $display("%b", result);

// TEST #620
// -914610.745122 + 0.000195807114372 = -914610.744926
// Expected Z = 11001001010111110100101100101100
#10 a = 32'b11001001010111110100101100101100; b = 32'b00111001010011010101000110010010; operation = 1'b0; $display("%b", result);

// TEST #621
// -396112.348733 - -0.000531825947132 = -396112.348201
// Expected Z = 11001000110000010110101000001011
#10 a = 32'b11001000110000010110101000001011; b = 32'b10111010000010110110101000111100; operation = 1'b1; $display("%b", result);

// TEST #622
// 863797.372273 - -0.000544625870979 = 863797.372817
// Expected Z = 01001001010100101110001101010110
#10 a = 32'b01001001010100101110001101010110; b = 32'b10111010000011101100010100111001; operation = 1'b1; $display("%b", result);

// TEST #623
// -934245.567588 + 0.000481650737117 = -934245.567106
// Expected Z = 11001001011001000001011001011001
#10 a = 32'b11001001011001000001011001011001; b = 32'b00111001111111001000011000010001; operation = 1'b0; $display("%b", result);

// TEST #624
// -308584.369761 + -0.000868423165281 = -308584.370629
// Expected Z = 11001000100101101010110100001100
#10 a = 32'b11001000100101101010110100001100; b = 32'b10111010011000111010011011100100; operation = 1'b0; $display("%b", result);

// TEST #625
// -691272.209142 + 0.000321831521696 = -691272.20882
// Expected Z = 11001001001010001100010010000011
#10 a = 32'b11001001001010001100010010000011; b = 32'b00111001101010001011101101111111; operation = 1'b0; $display("%b", result);

// TEST #626
// 652164.392943 - 1.36638388761e-05 = 652164.392929
// Expected Z = 01001001000111110011100001000110
#10 a = 32'b01001001000111110011100001000110; b = 32'b00110111011001010011110110111110; operation = 1'b1; $display("%b", result);

// TEST #627
// -81423.6669473 + -0.00024100034624 = -81423.6671883
// Expected Z = 11000111100111110000011111010101
#10 a = 32'b11000111100111110000011111010101; b = 32'b10111001011111001011010100001010; operation = 1'b0; $display("%b", result);

// TEST #628
// -348398.124946 + 0.000387035983353 = -348398.124559
// Expected Z = 11001000101010100001110111000100
#10 a = 32'b11001000101010100001110111000100; b = 32'b00111001110010101110101100010111; operation = 1'b0; $display("%b", result);

// TEST #629
// 911984.946244 + 0.000363855242641 = 911984.946608
// Expected Z = 01001001010111101010011100001111
#10 a = 32'b01001001010111101010011100001111; b = 32'b00111001101111101100001111010011; operation = 1'b0; $display("%b", result);

// TEST #630
// 753940.918055 + -0.000990842648094 = 753940.917064
// Expected Z = 01001001001110000001000101001111
#10 a = 32'b01001001001110000001000101001111; b = 32'b10111010100000011101111100101010; operation = 1'b0; $display("%b", result);

// TEST #631
// 92614.962438 + -0.000509670769691 = 92614.9619283
// Expected Z = 01000111101101001110001101111011
#10 a = 32'b01000111101101001110001101111011; b = 32'b10111010000001011001101101101101; operation = 1'b0; $display("%b", result);

// TEST #632
// 440881.010505 - -0.000202644600211 = 440881.010708
// Expected Z = 01001000110101110100011000100000
#10 a = 32'b01001000110101110100011000100000; b = 32'b10111001010101000111110011111111; operation = 1'b1; $display("%b", result);

// TEST #633
// 141409.278143 + 0.000974876191007 = 141409.279117
// Expected Z = 01001000000010100001100001010010
#10 a = 32'b01001000000010100001100001010010; b = 32'b00111010011111111000111011010101; operation = 1'b0; $display("%b", result);

// TEST #634
// -795870.354364 - 0.000516682031072 = -795870.35488
// Expected Z = 11001001010000100100110111100110
#10 a = 32'b11001001010000100100110111100110; b = 32'b00111010000001110111000111110010; operation = 1'b1; $display("%b", result);

// TEST #635
// 737126.174333 - -0.000402481045886 = 737126.174735
// Expected Z = 01001001001100111111011001100011
#10 a = 32'b01001001001100111111011001100011; b = 32'b10111001110100110000010000010111; operation = 1'b1; $display("%b", result);

// TEST #636
// -767616.292543 - 0.000965070798528 = -767616.293508
// Expected Z = 11001001001110110110100000000101
#10 a = 32'b11001001001110110110100000000101; b = 32'b00111010011111001111110011001110; operation = 1'b1; $display("%b", result);

// TEST #637
// -929057.050128 - 0.000317307250346 = -929057.050446
// Expected Z = 11001001011000101101001000010001
#10 a = 32'b11001001011000101101001000010001; b = 32'b00111001101001100101110001000010; operation = 1'b1; $display("%b", result);

// TEST #638
// -914490.912937 - 0.000384121955335 = -914490.913321
// Expected Z = 11001001010111110100001110101111
#10 a = 32'b11001001010111110100001110101111; b = 32'b00111001110010010110001111111010; operation = 1'b1; $display("%b", result);

// TEST #639
// 290164.101779 + -0.000123733450662 = 290164.101655
// Expected Z = 01001000100011011010111010000011
#10 a = 32'b01001000100011011010111010000011; b = 32'b10111001000000011011111001110010; operation = 1'b0; $display("%b", result);

// TEST #640
// -516708.592947 + 0.000600107471492 = -516708.592347
// Expected Z = 11001000111111000100110010010011
#10 a = 32'b11001000111111000100110010010011; b = 32'b00111010000111010101000010001000; operation = 1'b0; $display("%b", result);

// TEST #641
// -190455.699984 + -0.000768374817702 = -190455.700752
// Expected Z = 11001000001110011111110111101101
#10 a = 32'b11001000001110011111110111101101; b = 32'b10111010010010010110110011000011; operation = 1'b0; $display("%b", result);

// TEST #642
// 904573.766026 - 0.000281369600233 = 904573.765745
// Expected Z = 01001001010111001101011111011100
#10 a = 32'b01001001010111001101011111011100; b = 32'b00111001100100111000010011001010; operation = 1'b1; $display("%b", result);

// TEST #643
// -402898.222341 + -0.000410465423228 = -402898.222751
// Expected Z = 11001000110001001011101001000111
#10 a = 32'b11001000110001001011101001000111; b = 32'b10111001110101110011001110111101; operation = 1'b0; $display("%b", result);

// TEST #644
// 169214.745168 + -0.000313035115748 = 169214.744855
// Expected Z = 01001000001001010011111110110000
#10 a = 32'b01001000001001010011111110110000; b = 32'b10111001101001000001111011011101; operation = 1'b0; $display("%b", result);

// TEST #645
// 635340.80838 + 0.000522395872613 = 635340.808903
// Expected Z = 01001001000110110001110011001101
#10 a = 32'b01001001000110110001110011001101; b = 32'b00111010000010001111000101100101; operation = 1'b0; $display("%b", result);

// TEST #646
// -859052.267901 + -0.000565668513049 = -859052.268467
// Expected Z = 11001001010100011011101011000100
#10 a = 32'b11001001010100011011101011000100; b = 32'b10111010000101000100100101011111; operation = 1'b0; $display("%b", result);

// TEST #647
// -259187.03276 + -0.000237273847004 = -259187.032997
// Expected Z = 11001000011111010001110011000010
#10 a = 32'b11001000011111010001110011000010; b = 32'b10111001011110001100110010110111; operation = 1'b0; $display("%b", result);

// TEST #648
// -346440.97029 - -0.000676877709938 = -346440.969613
// Expected Z = 11001000101010010010100100011111
#10 a = 32'b11001000101010010010100100011111; b = 32'b10111010001100010111000001111111; operation = 1'b1; $display("%b", result);

// TEST #649
// -515888.104134 + -0.000547857100335 = -515888.104682
// Expected Z = 11001000111110111110011000000011
#10 a = 32'b11001000111110111110011000000011; b = 32'b10111010000011111001111000010001; operation = 1'b0; $display("%b", result);

// TEST #650
// 475101.443502 + 0.00075340853479 = 475101.444255
// Expected Z = 01001000111001111111101110101110
#10 a = 32'b01001000111001111111101110101110; b = 32'b00111010010001011000000001100100; operation = 1'b0; $display("%b", result);

// TEST #651
// 119293.647871 - -0.000886422796865 = 119293.648758
// Expected Z = 01000111111010001111111011010011
#10 a = 32'b01000111111010001111111011010011; b = 32'b10111010011010000101111011010100; operation = 1'b1; $display("%b", result);

// TEST #652
// 135098.520851 - -7.785931579e-05 = 135098.520928
// Expected Z = 01001000000000111110111010100001
#10 a = 32'b01001000000000111110111010100001; b = 32'b10111000101000110100100001100111; operation = 1'b1; $display("%b", result);

// TEST #653
// -92398.9404085 - -2.61225053947e-06 = -92398.9404059
// Expected Z = 11000111101101000111011101111000
#10 a = 32'b11000111101101000111011101111000; b = 32'b10110110001011110100111000011111; operation = 1'b1; $display("%b", result);

// TEST #654
// 427396.085508 - 0.000669707711332 = 427396.084838
// Expected Z = 01001000110100001011000010000011
#10 a = 32'b01001000110100001011000010000011; b = 32'b00111010001011111000111101010011; operation = 1'b1; $display("%b", result);

// TEST #655
// 256102.396709 + 0.000738783867066 = 256102.397447
// Expected Z = 01001000011110100001100110011001
#10 a = 32'b01001000011110100001100110011001; b = 32'b00111010010000011010101011110010; operation = 1'b0; $display("%b", result);

// TEST #656
// 714915.362463 + 0.000627513408087 = 714915.363091
// Expected Z = 01001001001011101000101000110110
#10 a = 32'b01001001001011101000101000110110; b = 32'b00111010001001000111111110110110; operation = 1'b0; $display("%b", result);

// TEST #657
// 12795.4730208 - -0.000994715691474 = 12795.4740155
// Expected Z = 01000110010001111110110111100101
#10 a = 32'b01000110010001111110110111100100; b = 32'b10111010100000100110000100011111; operation = 1'b1; $display("%b", result);

// TEST #658
// -294180.875482 - -0.000734333020665 = -294180.874748
// Expected Z = 11001000100011111010010010011100
#10 a = 32'b11001000100011111010010010011100; b = 32'b10111010010000001000000001000001; operation = 1'b1; $display("%b", result);

// TEST #659
// 591244.114971 + -0.000823385815704 = 591244.114148
// Expected Z = 01001001000100000101100011000010
#10 a = 32'b01001001000100000101100011000010; b = 32'b10111010010101111101100001111101; operation = 1'b0; $display("%b", result);

// TEST #660
// 233092.287186 - 5.92125158641e-05 = 233092.287127
// Expected Z = 01001000011000111010000100010010
#10 a = 32'b01001000011000111010000100010010; b = 32'b00111000011110000101101011110100; operation = 1'b1; $display("%b", result);

// TEST #661
// 796663.461968 - -8.07386085476e-05 = 796663.462049
// Expected Z = 01001001010000100111111101110111
#10 a = 32'b01001001010000100111111101110111; b = 32'b10111000101010010101001000110110; operation = 1'b1; $display("%b", result);

// TEST #662
// 917977.868522 - 0.000927904236882 = 917977.867594
// Expected Z = 01001001011000000001110110011110
#10 a = 32'b01001001011000000001110110011110; b = 32'b00111010011100110011111010011001; operation = 1'b1; $display("%b", result);

// TEST #663
// -751575.039906 - 0.000590219392366 = -751575.040496
// Expected Z = 11001001001101110111110101110001
#10 a = 32'b11001001001101110111110101110001; b = 32'b00111010000110101011100011110100; operation = 1'b1; $display("%b", result);

// TEST #664
// -413243.470218 - -0.00031261863242 = -413243.469905
// Expected Z = 11001000110010011100011101101111
#10 a = 32'b11001000110010011100011101101111; b = 32'b10111001101000111110011011110110; operation = 1'b1; $display("%b", result);

// TEST #665
// -116492.9647 - -6.22351573672e-05 = -116492.964638
// Expected Z = 11000111111000111000011001111011
#10 a = 32'b11000111111000111000011001111011; b = 32'b10111000100000101000010000111111; operation = 1'b1; $display("%b", result);

// TEST #666
// 876429.984053 - 0.00014574628045 = 876429.983907
// Expected Z = 01001001010101011111100011100000
#10 a = 32'b01001001010101011111100011100000; b = 32'b00111001000110001101001101111000; operation = 1'b1; $display("%b", result);

// TEST #667
// 766512.79207 - -0.00023132516745 = 766512.792301
// Expected Z = 01001001001110110010001100001101
#10 a = 32'b01001001001110110010001100001101; b = 32'b10111001011100101000111111100000; operation = 1'b1; $display("%b", result);

// TEST #668
// -553938.853336 - 0.000548591213821 = -553938.853885
// Expected Z = 11001001000001110011110100101110
#10 a = 32'b11001001000001110011110100101110; b = 32'b00111010000011111100111101010101; operation = 1'b1; $display("%b", result);

// TEST #669
// -666706.249696 - 0.000338889375355 = -666706.250035
// Expected Z = 11001001001000101100010100100100
#10 a = 32'b11001001001000101100010100100100; b = 32'b00111001101100011010110011110110; operation = 1'b1; $display("%b", result);

// TEST #670
// 371233.317583 - 0.00085327723152 = 371233.31673
// Expected Z = 01001000101101010100010000101010
#10 a = 32'b01001000101101010100010000101010; b = 32'b00111010010111111010111001110111; operation = 1'b1; $display("%b", result);

// TEST #671
// -150777.142839 - -0.000446479284804 = -150777.142392
// Expected Z = 11001000000100110011111001001001
#10 a = 32'b11001000000100110011111001001001; b = 32'b10111001111010100001010101101111; operation = 1'b1; $display("%b", result);

// TEST #672
// -438456.038269 + 0.000105196320263 = -438456.038164
// Expected Z = 11001000110101100001011100000001
#10 a = 32'b11001000110101100001011100000001; b = 32'b00111000110111001001110011011000; operation = 1'b0; $display("%b", result);

// TEST #673
// -250883.627804 - 0.000484784684931 = -250883.628289
// Expected Z = 11001000011101010000000011101000
#10 a = 32'b11001000011101010000000011101000; b = 32'b00111001111111100010101010110011; operation = 1'b1; $display("%b", result);

// TEST #674
// -770806.307141 + 0.000148534136392 = -770806.306992
// Expected Z = 11001001001111000010111101100101
#10 a = 32'b11001001001111000010111101100101; b = 32'b00111001000110111011111111010100; operation = 1'b0; $display("%b", result);

// TEST #675
// 597860.088808 + -0.000274097157769 = 597860.088534
// Expected Z = 01001001000100011111011001000001
#10 a = 32'b01001001000100011111011001000001; b = 32'b10111001100011111011010010110011; operation = 1'b0; $display("%b", result);

// TEST #676
// -165299.002691 + -0.000812193776111 = -165299.003503
// Expected Z = 11001000001000010110110011000000
#10 a = 32'b11001000001000010110110011000000; b = 32'b10111010010101001110100101100111; operation = 1'b0; $display("%b", result);

// TEST #677
// 255513.216674 + 0.000652558616588 = 255513.217327
// Expected Z = 01001000011110011000011001001110
#10 a = 32'b01001000011110011000011001001110; b = 32'b00111010001010110001000001111000; operation = 1'b0; $display("%b", result);

// TEST #678
// 830742.535347 + 8.89353378636e-05 = 830742.535436
// Expected Z = 01001001010010101101000101101001
#10 a = 32'b01001001010010101101000101101001; b = 32'b00111000101110101000001011001100; operation = 1'b0; $display("%b", result);

// TEST #679
// 657437.377445 - -0.000201833115906 = 657437.377647
// Expected Z = 01001001001000001000000111010110
#10 a = 32'b01001001001000001000000111010110; b = 32'b10111001010100111010001100101010; operation = 1'b1; $display("%b", result);

// TEST #680
// -294025.739096 + 0.000806874804834 = -294025.73829
// Expected Z = 11001000100011111001000100111000
#10 a = 32'b11001000100011111001000100111000; b = 32'b00111010010100111000010001110100; operation = 1'b0; $display("%b", result);

// TEST #681
// 303666.389122 - -0.000565189861746 = 303666.389687
// Expected Z = 01001000100101000100011001001100
#10 a = 32'b01001000100101000100011001001100; b = 32'b10111010000101000010100101000000; operation = 1'b1; $display("%b", result);

// TEST #682
// 984389.020918 - 0.000494031759972 = 984389.020424
// Expected Z = 01001001011100000101010001010000
#10 a = 32'b01001001011100000101010001010000; b = 32'b00111010000000011000000111101001; operation = 1'b1; $display("%b", result);

// TEST #683
// 506566.864365 + -0.000428869310005 = 506566.863936
// Expected Z = 01001000111101110101100011011100
#10 a = 32'b01001000111101110101100011011100; b = 32'b10111001111000001101100111011101; operation = 1'b0; $display("%b", result);

// TEST #684
// 454174.748986 - -0.000123164866499 = 454174.749109
// Expected Z = 01001000110111011100001111011000
#10 a = 32'b01001000110111011100001111011000; b = 32'b10111001000000010010010111010001; operation = 1'b1; $display("%b", result);

// TEST #685
// 929084.068876 + 0.000547135576715 = 929084.069423
// Expected Z = 01001001011000101101001111000001
#10 a = 32'b01001001011000101101001111000001; b = 32'b00111010000011110110110110100110; operation = 1'b0; $display("%b", result);

// TEST #686
// -189907.706849 - -0.000217568936685 = -189907.706631
// Expected Z = 11001000001110010111010011101101
#10 a = 32'b11001000001110010111010011101101; b = 32'b10111001011001000010001100110111; operation = 1'b1; $display("%b", result);

// TEST #687
// 901474.73692 - -0.000438418652136 = 901474.737358
// Expected Z = 01001001010111000001011000101100
#10 a = 32'b01001001010111000001011000101100; b = 32'b10111001111001011101101110001110; operation = 1'b1; $display("%b", result);

// TEST #688
// 28784.8262888 + 0.000347745322157 = 28784.8266366
// Expected Z = 01000110111000001110000110100111
#10 a = 32'b01000110111000001110000110100111; b = 32'b00111001101101100101000110010110; operation = 1'b0; $display("%b", result);

// TEST #689
// -551920.527443 + -0.000211708591429 = -551920.527655
// Expected Z = 11001001000001101011111100001000
#10 a = 32'b11001001000001101011111100001000; b = 32'b10111001010111011111111000011000; operation = 1'b0; $display("%b", result);

// TEST #690
// -792532.236687 - -0.000907373880276 = -792532.235779
// Expected Z = 11001001010000010111110101000100
#10 a = 32'b11001001010000010111110101000100; b = 32'b10111010011011011101110011010101; operation = 1'b1; $display("%b", result);

// TEST #691
// -146099.662966 - 0.00062615399408 = -146099.663592
// Expected Z = 11001000000011101010110011101010
#10 a = 32'b11001000000011101010110011101010; b = 32'b00111010001001000010010001111100; operation = 1'b1; $display("%b", result);

// TEST #692
// 993240.719887 - 0.000261106531406 = 993240.719626
// Expected Z = 01001001011100100111110110001100
#10 a = 32'b01001001011100100111110110001100; b = 32'b00111001100010001110010100100000; operation = 1'b1; $display("%b", result);

// TEST #693
// 703737.395803 - -0.000119831842525 = 703737.395923
// Expected Z = 01001001001010111100111110010110
#10 a = 32'b01001001001010111100111110010110; b = 32'b10111000111110110100111000111011; operation = 1'b1; $display("%b", result);

// TEST #694
// 371636.705418 + -0.000594410341839 = 371636.704824
// Expected Z = 01001000101101010111011010010111
#10 a = 32'b01001000101101010111011010010111; b = 32'b10111010000110111101001000110100; operation = 1'b0; $display("%b", result);

// TEST #695
// -999701.053476 + 0.000262754916062 = -999701.053213
// Expected Z = 11001001011101000001000101010001
#10 a = 32'b11001001011101000001000101010001; b = 32'b00111001100010011100001001011110; operation = 1'b0; $display("%b", result);

// TEST #696
// 668019.047268 + -0.000329962251131 = 668019.046938
// Expected Z = 01001001001000110001011100110001
#10 a = 32'b01001001001000110001011100110001; b = 32'b10111001101011001111111011001001; operation = 1'b0; $display("%b", result);

// TEST #697
// -213909.823353 + -0.000199824062767 = -213909.823553
// Expected Z = 11001000010100001110010101110101
#10 a = 32'b11001000010100001110010101110101; b = 32'b10111001010100011000011111011101; operation = 1'b0; $display("%b", result);

// TEST #698
// 140161.521586 - -0.000602700187201 = 140161.522189
// Expected Z = 01001000000010001110000001100001
#10 a = 32'b01001000000010001110000001100001; b = 32'b10111010000111011111111010000110; operation = 1'b1; $display("%b", result);

// TEST #699
// 831525.267422 + -0.000847007742641 = 831525.266575
// Expected Z = 01001001010010110000001001010100
#10 a = 32'b01001001010010110000001001010100; b = 32'b10111010010111100000100110111010; operation = 1'b0; $display("%b", result);

// TEST #700
// -431942.787899 + -0.000235486628418 = -431942.788135
// Expected Z = 11001000110100101110100011011001
#10 a = 32'b11001000110100101110100011011001; b = 32'b10111001011101101110110011110110; operation = 1'b0; $display("%b", result);

// TEST #701
// 0.872279998182 - -0.00069284770941 = 0.872972845891
// Expected Z = 00111111010111110111101100100110
#10 a = 32'b00111111010111110100110110111110; b = 32'b10111010001101011010000000111001; operation = 1'b1; $display("%b", result);

// TEST #702
// 0.662905845654 - 0.000223495891483 = 0.662682349762
// Expected Z = 00111111001010011010010110001101
#10 a = 32'b00111111001010011011010000110011; b = 32'b00111001011010100101101000111001; operation = 1'b1; $display("%b", result);

// TEST #703
// 0.340791571618 + 0.000945056896973 = 0.341736628515
// Expected Z = 00111110101011101111100000011010
#10 a = 32'b00111110101011100111110000111100; b = 32'b00111010011101111011110110110010; operation = 1'b0; $display("%b", result);

// TEST #704
// -0.823463554519 - -0.000318256339988 = -0.823145298179
// Expected Z = 10111111010100101011100110100110
#10 a = 32'b10111111010100101100111010000010; b = 32'b10111001101001101101101110100101; operation = 1'b1; $display("%b", result);

// TEST #705
// -0.775036157732 - -0.00069416369011 = -0.774341994042
// Expected Z = 10111111010001100011101101000111
#10 a = 32'b10111111010001100110100011000101; b = 32'b10111010001101011111100010001001; operation = 1'b1; $display("%b", result);

// TEST #706
// 0.662286742394 - -0.000517367815331 = 0.662804110209
// Expected Z = 00111111001010011010110110001000
#10 a = 32'b00111111001010011000101110100000; b = 32'b10111010000001111001111111110111; operation = 1'b1; $display("%b", result);

// TEST #707
// 0.0128880632498 + -3.89797329293e-05 = 0.0128490835168
// Expected Z = 00111100010100101000010011110110
#10 a = 32'b00111100010100110010100001110101; b = 32'b10111000001000110111111000101011; operation = 1'b0; $display("%b", result);

// TEST #708
// 0.432475033113 + -0.000986947665789 = 0.431488085447
// Expected Z = 00111110110111001110110000000010
#10 a = 32'b00111110110111010110110101011110; b = 32'b10111010100000010101110001111000; operation = 1'b0; $display("%b", result);

// TEST #709
// 0.972217987169 - -0.000996498089077 = 0.973214485258
// Expected Z = 00111111011110010010010010010110
#10 a = 32'b00111111011110001110001101000111; b = 32'b10111010100000101001110011101101; operation = 1'b1; $display("%b", result);

// TEST #710
// 0.168106458889 + 9.40083514231e-05 = 0.168200467241
// Expected Z = 00111110001011000011110010111110
#10 a = 32'b00111110001011000010010000011001; b = 32'b00111000110001010010011001011001; operation = 1'b0; $display("%b", result);

// TEST #711
// -0.308574970359 + -0.000948162339307 = -0.309523132698
// Expected Z = 10111110100111100111100111010001
#10 a = 32'b10111110100111011111110110001010; b = 32'b10111010011110001000111000011001; operation = 1'b0; $display("%b", result);

// TEST #712
// 0.737514380465 + -0.000520266381139 = 0.736994114083
// Expected Z = 00111111001111001010101110100101
#10 a = 32'b00111111001111001100110110111110; b = 32'b10111010000010000110001001111100; operation = 1'b0; $display("%b", result);

// TEST #713
// -0.943603107538 + 0.000226852439215 = -0.943376255099
// Expected Z = 10111111011100011000000100011011
#10 a = 32'b10111111011100011000111111111001; b = 32'b00111001011011011101111100111101; operation = 1'b0; $display("%b", result);

// TEST #714
// -0.768522894947 - -0.000338153991897 = -0.768184740955
// Expected Z = 10111111010001001010011111000001
#10 a = 32'b10111111010001001011110111101011; b = 32'b10111001101100010100101001000011; operation = 1'b1; $display("%b", result);

// TEST #715
// -0.11433562944 - 0.000437318876895 = -0.114772948316
// Expected Z = 10111101111010110000111000010100
#10 a = 32'b10111101111010100010100011001100; b = 32'b00111001111001010100011111110010; operation = 1'b1; $display("%b", result);

// TEST #716
// -0.473533349194 + 0.000152461601719 = -0.473380887592
// Expected Z = 10111110111100100101111011111011
#10 a = 32'b10111110111100100111001011110111; b = 32'b00111001000111111101111000011001; operation = 1'b0; $display("%b", result);

// TEST #717
// 0.63114777628 + -0.000677730726036 = 0.630470045553
// Expected Z = 00111111001000010110011001111100
#10 a = 32'b00111111001000011001001011100111; b = 32'b10111010001100011010100110111101; operation = 1'b0; $display("%b", result);

// TEST #718
// 0.737484360935 + -2.29309154758e-05 = 0.73746143002
// Expected Z = 00111111001111001100101001000110
#10 a = 32'b00111111001111001100101111000110; b = 32'b10110111110000000101101111000100; operation = 1'b0; $display("%b", result);

// TEST #719
// 0.617611743362 + -0.000283094110644 = 0.617328649252
// Expected Z = 00111111000111100000100101000000
#10 a = 32'b00111111000111100001101111001110; b = 32'b10111001100101000110110001000000; operation = 1'b0; $display("%b", result);

// TEST #720
// 0.083765052033 - -0.000511472380664 = 0.0842765244137
// Expected Z = 00111101101011001001100100101100
#10 a = 32'b00111101101010111000110100000011; b = 32'b10111010000001100001010001010101; operation = 1'b1; $display("%b", result);

// TEST #721
// -0.553273436402 - -0.000167728678858 = -0.553105707723
// Expected Z = 10111111000011011001100001010110
#10 a = 32'b10111111000011011010001101010100; b = 32'b10111001001011111110000001010011; operation = 1'b1; $display("%b", result);

// TEST #722
// -0.228755585899 - -0.000926003635397 = -0.227829582264
// Expected Z = 10111110011010010100110000101000
#10 a = 32'b10111110011010100011111011101000; b = 32'b10111010011100101011111100001101; operation = 1'b1; $display("%b", result);

// TEST #723
// 0.83073075573 + -0.000506023308966 = 0.830224732421
// Expected Z = 00111111010101001000100110011100
#10 a = 32'b00111111010101001010101011000101; b = 32'b10111010000001001010011010100110; operation = 1'b0; $display("%b", result);

// TEST #724
// 0.674185323514 + -0.000157630959553 = 0.674027692554
// Expected Z = 00111111001011001000110100010100
#10 a = 32'b00111111001011001001011101101001; b = 32'b10111001001001010100100110111101; operation = 1'b0; $display("%b", result);

// TEST #725
// 0.312935772455 - 0.000612541086056 = 0.312323231369
// Expected Z = 00111110100111111110100011010101
#10 a = 32'b00111110101000000011100100011110; b = 32'b00111010001000001001001011110000; operation = 1'b1; $display("%b", result);

// TEST #726
// 0.412261547022 - -0.000824868879404 = 0.413086415901
// Expected Z = 00111110110100111000000000010000
#10 a = 32'b00111110110100110001001111110010; b = 32'b10111010010110000011110000000011; operation = 1'b1; $display("%b", result);

// TEST #727
// 0.411587120951 - 0.000393161681786 = 0.411193959269
// Expected Z = 00111110110100101000100000000100
#10 a = 32'b00111110110100101011101110001100; b = 32'b00111001110011100010000101000101; operation = 1'b1; $display("%b", result);

// TEST #728
// -0.163095765485 - -0.000975772242773 = -0.162119993242
// Expected Z = 10111110001001100000001011001001
#10 a = 32'b10111110001001110000001010010100; b = 32'b10111010011111111100101011110111; operation = 1'b1; $display("%b", result);

// TEST #729
// 0.842023177969 + -0.000241501084805 = 0.841781676884
// Expected Z = 00111111010101110111111100000001
#10 a = 32'b00111111010101111000111011010101; b = 32'b10111001011111010011101101110100; operation = 1'b0; $display("%b", result);

// TEST #730
// 0.666230299938 - 0.000173594463513 = 0.666056705475
// Expected Z = 00111111001010101000001010110001
#10 a = 32'b00111111001010101000111000010010; b = 32'b00111001001101100000011011101001; operation = 1'b1; $display("%b", result);

// TEST #731
// 1.97260125218e-05 + -0.000893246465021 = -0.000873520452499
// Expected Z = 10111010011001001111110011110111
#10 a = 32'b00110111101001010111100101001010; b = 32'b10111010011010100010100011000001; operation = 1'b0; $display("%b", result);

// TEST #732
// 0.11794773809 - -4.86696254974e-05 = 0.117996407715
// Expected Z = 00111101111100011010100000011010
#10 a = 32'b00111101111100011000111010010101; b = 32'b10111000010011000010001010011101; operation = 1'b1; $display("%b", result);

// TEST #733
// 0.535949103281 + 0.000671314841345 = 0.536620418122
// Expected Z = 00111111000010010101111111110101
#10 a = 32'b00111111000010010011001111110110; b = 32'b00111010001011111111101100101101; operation = 1'b0; $display("%b", result);

// TEST #734
// -0.564956252883 - -0.000442375515117 = -0.564513877368
// Expected Z = 10111111000100001000001111111011
#10 a = 32'b10111111000100001010000011111001; b = 32'b10111001111001111110111010100011; operation = 1'b1; $display("%b", result);

// TEST #735
// -0.285489022091 + 0.0002340100447 = -0.285255012047
// Expected Z = 10111110100100100000110011110010
#10 a = 32'b10111110100100100010101110011110; b = 32'b00111001011101010110000010011000; operation = 1'b0; $display("%b", result);

// TEST #736
// -0.553209743667 + -0.000955382655153 = -0.554165126322
// Expected Z = 10111111000011011101110111000100
#10 a = 32'b10111111000011011001111100100111; b = 32'b10111010011110100111001010100101; operation = 1'b0; $display("%b", result);

// TEST #737
// -0.184757587856 - -8.72527604163e-05 = -0.184670335096
// Expected Z = 10111110001111010001101000111000
#10 a = 32'b10111110001111010011000100011000; b = 32'b10111000101101101111101101111000; operation = 1'b1; $display("%b", result);

// TEST #738
// -0.518409197915 - -0.000630653787424 = -0.517778544127
// Expected Z = 10111111000001001000110100100010
#10 a = 32'b10111111000001001011011001110111; b = 32'b10111010001001010101001001110110; operation = 1'b1; $display("%b", result);

// TEST #739
// -0.194835052015 + -0.000181857029532 = -0.195016909044
// Expected Z = 10111110010001111011001010000011
#10 a = 32'b10111110010001111000001011010111; b = 32'b10111001001111101011000011100000; operation = 1'b0; $display("%b", result);

// TEST #740
// 0.513932275986 - 0.000247403286768 = 0.513684872699
// Expected Z = 00111111000000111000000011011010
#10 a = 32'b00111111000000111001000100010001; b = 32'b00111001100000011011010111101000; operation = 1'b1; $display("%b", result);

// TEST #741
// 0.349447203021 + -0.000728015792609 = 0.348719187228
// Expected Z = 00111110101100101000101101010010
#10 a = 32'b00111110101100101110101010111110; b = 32'b10111010001111101101100001010000; operation = 1'b0; $display("%b", result);

// TEST #742
// 0.419313153773 - 0.000417795447293 = 0.418895358326
// Expected Z = 00111110110101100111100101110100
#10 a = 32'b00111110110101101011000000110111; b = 32'b00111001110110110000101110001110; operation = 1'b1; $display("%b", result);

// TEST #743
// 0.149206978756 - -0.000767081489766 = 0.149974060245
// Expected Z = 00111110000110011001001011001101
#10 a = 32'b00111110000110001100100110110111; b = 32'b10111010010010010001010111111000; operation = 1'b1; $display("%b", result);

// TEST #744
// -0.543579995881 - -0.000822080598748 = -0.542757915282
// Expected Z = 10111111000010101111001000101111
#10 a = 32'b10111111000010110010100000001111; b = 32'b10111010010101111000000011100101; operation = 1'b1; $display("%b", result);

// TEST #745
// 0.368600818058 - -0.000254078898205 = 0.368854896956
// Expected Z = 00111110101111001101101010001101
#10 a = 32'b00111110101111001011100100111111; b = 32'b10111001100001010011010111100100; operation = 1'b1; $display("%b", result);

// TEST #746
// 0.82202483828 - -0.000288297021818 = 0.822313135302
// Expected Z = 00111111010100101000001100011101
#10 a = 32'b00111111010100100111000000111000; b = 32'b10111001100101110010011010010010; operation = 1'b1; $display("%b", result);

// TEST #747
// -0.412770819364 + -0.000465697687304 = -0.413236517051
// Expected Z = 10111110110100111001001110111101
#10 a = 32'b10111110110100110101011010110010; b = 32'b10111001111101000010100011100011; operation = 1'b0; $display("%b", result);

// TEST #748
// -0.31651302449 - -0.000424621170756 = -0.316088403319
// Expected Z = 10111110101000011101011001010111
#10 a = 32'b10111110101000100000110111111111; b = 32'b10111001110111101001111110110000; operation = 1'b1; $display("%b", result);

// TEST #749
// 0.369260698257 + 0.000964893681313 = 0.370225591938
// Expected Z = 00111110101111011000111000110101
#10 a = 32'b00111110101111010000111110111101; b = 32'b00111010011111001111000011101011; operation = 1'b0; $display("%b", result);

// TEST #750
// 0.481616962695 + -0.000348875608721 = 0.481268087086
// Expected Z = 00111110111101100110100011000101
#10 a = 32'b00111110111101101001011010000000; b = 32'b10111001101101101110100101001011; operation = 1'b0; $display("%b", result);

// TEST #751
// -0.559582325686 + 0.00077820928115 = -0.558804116405
// Expected Z = 10111111000011110000110111001001
#10 a = 32'b10111111000011110100000011001010; b = 32'b00111010010011000000000010111110; operation = 1'b0; $display("%b", result);

// TEST #752
// 0.0874591984426 - -0.000239607428297 = 0.0876988058709
// Expected Z = 00111101101100111001101101101110
#10 a = 32'b00111101101100110001110111001111; b = 32'b10111001011110110011111100100001; operation = 1'b1; $display("%b", result);

// TEST #753
// 0.737690587962 + -0.000819199174534 = 0.736871388787
// Expected Z = 00111111001111001010001110011010
#10 a = 32'b00111111001111001101100101001010; b = 32'b10111010010101101011111110000111; operation = 1'b0; $display("%b", result);

// TEST #754
// 0.0806524004958 + -1.69940186222e-05 = 0.0806354064772
// Expected Z = 00111101101001010010010000101101
#10 a = 32'b00111101101001010010110100010110; b = 32'b10110111100011101000111001100001; operation = 1'b0; $display("%b", result);

// TEST #755
// 0.885203353045 - -0.000309176897563 = 0.885512529943
// Expected Z = 00111111011000101011000011110011
#10 a = 32'b00111111011000101001110010110000; b = 32'b10111001101000100001100100000101; operation = 1'b1; $display("%b", result);

// TEST #756
// -0.658303849258 + -0.000398932411354 = -0.658702781669
// Expected Z = 10111111001010001010000010111111
#10 a = 32'b10111111001010001000011010011010; b = 32'b10111001110100010010011111001101; operation = 1'b0; $display("%b", result);

// TEST #757
// -0.40199717531 + -0.00069194919289 = -0.402689124503
// Expected Z = 10111110110011100010110101000101
#10 a = 32'b10111110110011011101001010010011; b = 32'b10111010001101010110001111101101; operation = 1'b0; $display("%b", result);

// TEST #758
// -0.284878942534 + 0.0004690087838 = -0.28440993375
// Expected Z = 10111110100100011001111000101110
#10 a = 32'b10111110100100011101101110100111; b = 32'b00111001111101011110010101001011; operation = 1'b0; $display("%b", result);

// TEST #759
// 0.178396918296 + -0.000668385255265 = 0.177728533041
// Expected Z = 00111110001101011111111001111000
#10 a = 32'b00111110001101101010110110101111; b = 32'b10111010001011110011011010010011; operation = 1'b0; $display("%b", result);

// TEST #760
// -0.155453865027 - -0.000644475637324 = -0.15480938939
// Expected Z = 10111110000111101000011001011010
#10 a = 32'b10111110000111110010111101001100; b = 32'b10111010001010001111001000000111; operation = 1'b1; $display("%b", result);

// TEST #761
// -0.223708869604 - -0.000472396363942 = -0.22323647324
// Expected Z = 10111110011001001001100000011010
#10 a = 32'b10111110011001010001001111110000; b = 32'b10111001111101111010101111110111; operation = 1'b1; $display("%b", result);

// TEST #762
// 0.337289323331 + 0.000364884192381 = 0.337654207523
// Expected Z = 00111110101011001110000100000011
#10 a = 32'b00111110101011001011000100110000; b = 32'b00111001101111110100110111101101; operation = 1'b0; $display("%b", result);

// TEST #763
// 0.997295269216 - -0.000938118024566 = 0.99823338724
// Expected Z = 00111111011111111000110000111001
#10 a = 32'b00111111011111110100111010111110; b = 32'b10111010011101011110110000001001; operation = 1'b1; $display("%b", result);

// TEST #764
// -0.535891380082 - 0.000666851269048 = -0.536558231351
// Expected Z = 10111111000010010101101111100001
#10 a = 32'b10111111000010010011000000101101; b = 32'b00111010001011101100111110100010; operation = 1'b1; $display("%b", result);

// TEST #765
// -0.818532573328 + 0.00031461819804 = -0.81821795513
// Expected Z = 10111111010100010111011010111011
#10 a = 32'b10111111010100011000101101011010; b = 32'b00111001101001001111001101010111; operation = 1'b0; $display("%b", result);

// TEST #766
// -0.129979280264 - 0.000299461642865 = -0.130278741907
// Expected Z = 10111110000001010110011111001010
#10 a = 32'b10111110000001010001100101001010; b = 32'b00111001100111010000000100010000; operation = 1'b1; $display("%b", result);

// TEST #767
// -0.964441233064 - 0.000986170788761 = -0.965427403853
// Expected Z = 10111111011101110010011001000000
#10 a = 32'b10111111011101101110010110011111; b = 32'b00111010100000010100001001100111; operation = 1'b1; $display("%b", result);

// TEST #768
// 0.302150789962 + -0.000533258479059 = 0.301617531483
// Expected Z = 00111110100110100110110110011101
#10 a = 32'b00111110100110101011001110000010; b = 32'b10111010000010111100101001011111; operation = 1'b0; $display("%b", result);

// TEST #769
// 0.251102663952 - 0.000444217557727 = 0.250658446394
// Expected Z = 00111110100000000101011001001110
#10 a = 32'b00111110100000001001000010000111; b = 32'b00111001111010001110010111011111; operation = 1'b1; $display("%b", result);

// TEST #770
// -0.747159473315 - -0.000382212706409 = -0.746777260608
// Expected Z = 10111111001111110010110011001011
#10 a = 32'b10111111001111110100010111011000; b = 32'b10111001110010000110001110111001; operation = 1'b1; $display("%b", result);

// TEST #771
// -0.0597062466439 - -0.000320315111252 = -0.0593859315327
// Expected Z = 10111101011100110011111010101010
#10 a = 32'b10111101011101001000111010001010; b = 32'b10111001101001111110111111110111; operation = 1'b1; $display("%b", result);

// TEST #772
// -0.469311794978 - 0.000813646332134 = -0.47012544131
// Expected Z = 10111110111100001011010001001000
#10 a = 32'b10111110111100000100100110100011; b = 32'b00111010010101010100101011100010; operation = 1'b1; $display("%b", result);

// TEST #773
// 0.330030150445 + 0.000870190303529 = 0.330900340749
// Expected Z = 00111110101010010110101111000101
#10 a = 32'b00111110101010001111100110110110; b = 32'b00111010011001000001110101111100; operation = 1'b0; $display("%b", result);

// TEST #774
// 0.993373299152 - 3.01489767906e-05 = 0.993343150175
// Expected Z = 00111111011111100100101110111101
#10 a = 32'b00111111011111100100110110110110; b = 32'b00110111111111001110100001101111; operation = 1'b1; $display("%b", result);

// TEST #775
// 0.878425673731 + 0.000287580700033 = 0.878713254431
// Expected Z = 00111111011000001111001101011010
#10 a = 32'b00111111011000001110000010000001; b = 32'b00111001100101101100011001101110; operation = 1'b0; $display("%b", result);

// TEST #776
// -0.781091184436 - -0.000489326613676 = -0.780601857823
// Expected Z = 10111111010001111101010110000110
#10 a = 32'b10111111010001111111010110011000; b = 32'b10111010000000000100011000100111; operation = 1'b1; $display("%b", result);

// TEST #777
// 0.486768601954 - -0.00075563876652 = 0.48752424072
// Expected Z = 00111110111110011001110011000111
#10 a = 32'b00111110111110010011100110111100; b = 32'b10111010010001100001011000001111; operation = 1'b1; $display("%b", result);

// TEST #778
// 0.122632479247 + -0.000792798167375 = 0.12183968108
// Expected Z = 00111101111110011000011100010101
#10 a = 32'b00111101111110110010011010111101; b = 32'b10111010010011111101001111001001; operation = 1'b0; $display("%b", result);

// TEST #779
// 0.0303651221956 + -2.12271681988e-05 = 0.0303438950274
// Expected Z = 00111100111110001001001111000011
#10 a = 32'b00111100111110001100000001000111; b = 32'b10110111101100100001000011111111; operation = 1'b0; $display("%b", result);

// TEST #780
// -0.798692779126 - -0.000493377782471 = -0.798199401343
// Expected Z = 10111111010011000101011011001100
#10 a = 32'b10111111010011000111011100100001; b = 32'b10111010000000010101011000000110; operation = 1'b1; $display("%b", result);

// TEST #781
// -0.726009011332 - -0.000955473997617 = -0.725053537334
// Expected Z = 10111111001110011001110100011100
#10 a = 32'b10111111001110011101101110111010; b = 32'b10111010011110100111100011000110; operation = 1'b1; $display("%b", result);

// TEST #782
// 0.760994273021 + 0.000923995803598 = 0.761918268825
// Expected Z = 00111111010000110000110100010011
#10 a = 32'b00111111010000101101000010000101; b = 32'b00111010011100100011100001001111; operation = 1'b0; $display("%b", result);

// TEST #783
// 0.783431967531 - 0.000545790669012 = 0.782886176862
// Expected Z = 00111111010010000110101100111010
#10 a = 32'b00111111010010001000111011111111; b = 32'b00111010000011110001001101100100; operation = 1'b1; $display("%b", result);

// TEST #784
// 0.855978557694 + 0.000575368039495 = 0.856553925734
// Expected Z = 00111111010110110100011100011110
#10 a = 32'b00111111010110110010000101101001; b = 32'b00111010000101101101010001001100; operation = 1'b0; $display("%b", result);

// TEST #785
// 0.897393341763 + -0.000523574533585 = 0.896869767229
// Expected Z = 00111111011001011001100101000010
#10 a = 32'b00111111011001011011101110010010; b = 32'b10111010000010010100000001111110; operation = 1'b0; $display("%b", result);

// TEST #786
// 0.32450936926 - 0.000419199974479 = 0.324090169285
// Expected Z = 00111110101001011110111100100110
#10 a = 32'b00111110101001100010011000011000; b = 32'b00111001110110111100100000010001; operation = 1'b1; $display("%b", result);

// TEST #787
// 0.691693391727 + 0.000468424921 = 0.692161816648
// Expected Z = 00111111001100010011000110000100
#10 a = 32'b00111111001100010001001011010001; b = 32'b00111001111101011001011011101110; operation = 1'b0; $display("%b", result);

// TEST #788
// -0.14296039649 - 0.000227160816148 = -0.143187557306
// Expected Z = 10111110000100101001111111000010
#10 a = 32'b10111110000100100110010000110110; b = 32'b00111001011011100011001000000100; operation = 1'b1; $display("%b", result);

// TEST #789
// -0.331994849862 - 0.000752086990818 = -0.332746936852
// Expected Z = 10111110101010100101110111001110
#10 a = 32'b10111110101010011111101100111011; b = 32'b00111010010001010010011110110100; operation = 1'b1; $display("%b", result);

// TEST #790
// 0.643995725069 - 0.000400220356319 = 0.643595504713
// Expected Z = 00111111001001001100001010101101
#10 a = 32'b00111111001001001101110011100111; b = 32'b00111001110100011101010010101011; operation = 1'b1; $display("%b", result);

// TEST #791
// 0.331229066979 + -0.000972825761583 = 0.330256241218
// Expected Z = 00111110101010010001011101011001
#10 a = 32'b00111110101010011001011011011011; b = 32'b10111010011111110000010100111011; operation = 1'b0; $display("%b", result);

// TEST #792
// -0.635249687794 + -0.000113414374888 = -0.635363102169
// Expected Z = 10111111001000101010011100101000
#10 a = 32'b10111111001000101001111110111001; b = 32'b10111000111011011101100011100001; operation = 1'b0; $display("%b", result);

// TEST #793
// -0.522037490167 - 0.000225957748361 = -0.522263447915
// Expected Z = 10111111000001011011001100001111
#10 a = 32'b10111111000001011010010001000000; b = 32'b00111001011011001110111100010010; operation = 1'b1; $display("%b", result);

// TEST #794
// 0.259568527244 - 0.000751539307566 = 0.258816987936
// Expected Z = 00111110100001001000001110101001
#10 a = 32'b00111110100001001110011000101010; b = 32'b00111010010001010000001011110011; operation = 1'b1; $display("%b", result);

// TEST #795
// -0.0872273782315 - -0.000542124403666 = -0.0866852538278
// Expected Z = 10111101101100011000100000001010
#10 a = 32'b10111101101100101010010001000101; b = 32'b10111010000011100001110101011010; operation = 1'b1; $display("%b", result);

// TEST #796
// 0.225453760735 - -0.000780880254233 = 0.22623464099
// Expected Z = 00111110011001111010101000001110
#10 a = 32'b00111110011001101101110101011010; b = 32'b10111010010011001011001111111101; operation = 1'b1; $display("%b", result);

// TEST #797
// -0.781678744819 - -0.000520671653998 = -0.781158073165
// Expected Z = 10111111010001111111100111111010
#10 a = 32'b10111111010010000001110000011001; b = 32'b10111010000010000111110110101111; operation = 1'b1; $display("%b", result);

// TEST #798
// -0.419180990929 - 0.000932359399102 = -0.420113350328
// Expected Z = 10111110110101110001100100011001
#10 a = 32'b10111110110101101001111011100100; b = 32'b00111010011101000110100110010101; operation = 1'b1; $display("%b", result);

// TEST #799
// -0.269910728223 + -0.000884878687515 = -0.27079560691
// Expected Z = 10111110100010101010010110111001
#10 a = 32'b10111110100010100011000110111101; b = 32'b10111010011001111111011100110100; operation = 1'b0; $display("%b", result);

// TEST #800
// -0.835916829353 - 0.000170180408025 = -0.836087009761
// Expected Z = 10111111010101100000100111001100
#10 a = 32'b10111111010101011111111010100101; b = 32'b00111001001100100111001001110101; operation = 1'b1; $display("%b", result);

// TEST #801
// 9.59372744104e-05 - 5.35351850464e-05 = 4.2402089364e-05
// Expected Z = 00111000001100011101100011100110
#10 a = 32'b00111000110010010011000111101111; b = 32'b00111000011000001000101011111000; operation = 1'b1; $display("%b", result);

// TEST #802
// -5.35918870683e-05 - -4.4126247365e-05 = -9.4656397033e-06
// Expected Z = 10110111000111101100111010011101
#10 a = 32'b10111000011000001100011111011010; b = 32'b10111000001110010001010000110011; operation = 1'b1; $display("%b", result);

// TEST #803
// 6.0591502736e-05 - -6.44405432517e-05 = 0.000125032045988
// Expected Z = 00111001000000110001101100001001
#10 a = 32'b00111000011111100010001110100001; b = 32'b10111000100001110010010001000001; operation = 1'b1; $display("%b", result);

// TEST #804
// -4.5872421152e-05 - -7.16475977529e-05 = 2.57751766009e-05
// Expected Z = 00110111110110000011011111000101
#10 a = 32'b10111000010000000110011100100011; b = 32'b10111000100101100100000110000011; operation = 1'b1; $display("%b", result);

// TEST #805
// 9.73636624943e-06 - 8.08271889053e-05 = -7.10908226559e-05
// Expected Z = 10111000100101010001011010011000
#10 a = 32'b00110111001000110101100101100000; b = 32'b00111000101010011000000111000100; operation = 1'b1; $display("%b", result);

// TEST #806
// -1.58985763901e-05 - -4.72026756101e-05 = 3.130409922e-05
// Expected Z = 00111000000000110100110010000101
#10 a = 32'b10110111100001010101110111101111; b = 32'b10111000010001011111101101111101; operation = 1'b1; $display("%b", result);

// TEST #807
// -6.58143147126e-05 + -2.36043919413e-05 = -8.94187066539e-05
// Expected Z = 10111000101110111000011001001101
#10 a = 32'b10111000100010100000010111001011; b = 32'b10110111110001100000001000001100; operation = 1'b0; $display("%b", result);

// TEST #808
// -6.91402444628e-05 + 8.28279207779e-06 = -6.0857452385e-05
// Expected Z = 10111000011111110100000100110001
#10 a = 32'b10111000100100001111111101100011; b = 32'b00110111000010101111011001010010; operation = 1'b0; $display("%b", result);

// TEST #809
// -4.89381640082e-05 - 8.28790371465e-05 = -0.000131817201155
// Expected Z = 10111001000010100011100001101001
#10 a = 32'b10111000010011010100001011110100; b = 32'b00111000101011011100111101011000; operation = 1'b1; $display("%b", result);

// TEST #810
// 4.24074025272e-05 + 5.26039178653e-05 = 9.50113203925e-05
// Expected Z = 00111000110001110100000011010000
#10 a = 32'b00111000001100011101111010011010; b = 32'b00111000010111001010001100000111; operation = 1'b0; $display("%b", result);

// TEST #811
// 1.33141571404e-05 + 2.89879571264e-05 = 4.23021142667e-05
// Expected Z = 00111000001100010110110110001101
#10 a = 32'b00110111010111110101111111011111; b = 32'b00110111111100110010101100101010; operation = 1'b0; $display("%b", result);

// TEST #812
// -7.34819444849e-06 - 3.07712594464e-05 = -3.81194538948e-05
// Expected Z = 10111000000111111110001001110100
#10 a = 32'b10110110111101101001000010000010; b = 32'b00111000000000010001000001100011; operation = 1'b1; $display("%b", result);

// TEST #813
// -6.10950332121e-06 + 4.97672823582e-05 = 4.3657779037e-05
// Expected Z = 00111000001101110001110100101111
#10 a = 32'b10110110110011010000000000111100; b = 32'b00111000010100001011110100110110; operation = 1'b0; $display("%b", result);

// TEST #814
// 3.88029552298e-06 + -2.33840675192e-05 = -1.95037719962e-05
// Expected Z = 10110111101000111001110000001000
#10 a = 32'b00110110100000100011001101111100; b = 32'b10110111110001000010100011100111; operation = 1'b0; $display("%b", result);

// TEST #815
// 8.25438582227e-05 - -6.48400761419e-05 = 0.000147383934365
// Expected Z = 00111001000110101000101100010011
#10 a = 32'b00111000101011010001101101100101; b = 32'b10111000100001111111101011000000; operation = 1'b1; $display("%b", result);

// TEST #816
// 7.52665857711e-06 + -4.33131369348e-05 = -3.57864783577e-05
// Expected Z = 10111000000101100001100101110000
#10 a = 32'b00110110111111001000110110000001; b = 32'b10111000001101011010101100100000; operation = 1'b0; $display("%b", result);

// TEST #817
// -9.97216025414e-05 + -7.29442478019e-05 = -0.000172665850343
// Expected Z = 10111001001101010000110110100011
#10 a = 32'b10111000110100010010000110100001; b = 32'b10111000100110001111100110100101; operation = 1'b0; $display("%b", result);

// TEST #818
// 9.63838581436e-05 + 8.83108448183e-05 = 0.000184694702962
// Expected Z = 00111001010000011010101010011011
#10 a = 32'b00111000110010100010000110110001; b = 32'b00111000101110010011001110000110; operation = 1'b0; $display("%b", result);

// TEST #819
// -4.04824177365e-05 - 5.3624211202e-05 = -9.41066289385e-05
// Expected Z = 10111000110001010101101100011101
#10 a = 32'b10111000001010011100101110101010; b = 32'b00111000011000001110101010001111; operation = 1'b1; $display("%b", result);

// TEST #820
// 8.59699652705e-05 + -5.44658605696e-05 = 3.15041047009e-05
// Expected Z = 00111000000001000010001101000110
#10 a = 32'b00111000101101000100101011000110; b = 32'b10111000011001000111001001000110; operation = 1'b0; $display("%b", result);

// TEST #821
// -2.67133212992e-06 - -2.70910648899e-05 = 2.441973276e-05
// Expected Z = 00110111110011001101100011111010
#10 a = 32'b10110110001100110100010100100011; b = 32'b10110111111000110100000110011110; operation = 1'b1; $display("%b", result);

// TEST #822
// -7.53127534808e-05 + -8.89209621719e-05 = -0.000164233715653
// Expected Z = 10111001001011000011011000100111
#10 a = 32'b10111000100111011111000100111010; b = 32'b10111000101110100111101100010100; operation = 1'b0; $display("%b", result);

// TEST #823
// -8.97623015595e-05 - -4.41077094417e-05 = -4.56545921178e-05
// Expected Z = 10111000001111110111110100111111
#10 a = 32'b10111000101111000011111011000101; b = 32'b10111000001110010000000001001011; operation = 1'b1; $display("%b", result);

// TEST #824
// -7.34679019132e-05 - 6.97030027817e-05 = -0.000143170904695
// Expected Z = 10111001000101100010000000100110
#10 a = 32'b10111000100110100001001011001000; b = 32'b00111000100100100010110110000100; operation = 1'b1; $display("%b", result);

// TEST #825
// -2.95600310034e-05 - -2.19940319383e-05 = -7.56599906517e-06
// Expected Z = 10110110111111011101111101110000
#10 a = 32'b10110111111101111111011110101111; b = 32'b10110111101110000111111111010011; operation = 1'b1; $display("%b", result);

// TEST #826
// 4.17309195378e-05 - -5.99765663185e-05 = 0.000101707485856
// Expected Z = 00111000110101010100101111001010
#10 a = 32'b00111000001011110000100000111100; b = 32'b10111000011110111000111101011001; operation = 1'b1; $display("%b", result);

// TEST #827
// 2.61034322125e-07 - 6.19416706661e-05 = -6.1680636344e-05
// Expected Z = 10111000100000010101101010001010
#10 a = 32'b00110100100011000010010001001001; b = 32'b00111000100000011110011010101110; operation = 1'b1; $display("%b", result);

// TEST #828
// 3.56433424099e-05 + -4.01044475722e-05 = -4.4611051623e-06
// Expected Z = 10110110100101011011000010011010
#10 a = 32'b00111000000101010111111110111111; b = 32'b10111000001010000011010111010011; operation = 1'b0; $display("%b", result);

// TEST #829
// -4.47112050543e-05 - 1.22546452413e-05 = -5.69658502956e-05
// Expected Z = 10111000011011101110111010011110
#10 a = 32'b10111000001110111000100001001010; b = 32'b00110111010011011001100101001101; operation = 1'b1; $display("%b", result);

// TEST #830
// -1.73430296936e-06 - -6.08430723532e-05 = 5.91087693839e-05
// Expected Z = 00111000011101111110101110001111
#10 a = 32'b10110101111010001100011000110010; b = 32'b10111000011111110011000111000000; operation = 1'b1; $display("%b", result);

// TEST #831
// 5.00438408039e-05 - -2.91897964433e-05 = 7.92336372472e-05
// Expected Z = 00111000101001100010101000111100
#10 a = 32'b00111000010100011110011000101010; b = 32'b10110111111101001101110010011100; operation = 1'b1; $display("%b", result);

// TEST #832
// -1.04241618225e-05 - -9.92160309694e-05 = 8.87918691469e-05
// Expected Z = 00111000101110100011010111000110
#10 a = 32'b10110111001011101110001101101111; b = 32'b10111000110100000001001000110011; operation = 1'b1; $display("%b", result);

// TEST #833
// -6.98324512912e-05 - -2.42050738883e-05 = -4.56273774028e-05
// Expected Z = 10111000001111110110000000000110
#10 a = 32'b10111000100100100111001100000011; b = 32'b10110111110010110000110000000000; operation = 1'b1; $display("%b", result);

// TEST #834
// -1.47878320882e-05 - -1.99853835965e-05 = 5.19755150826e-06
// Expected Z = 00110110101011100110011010100001
#10 a = 32'b10110111011110000001100101000001; b = 32'b10110111101001111010011001001001; operation = 1'b1; $display("%b", result);

// TEST #835
// 4.77182988816e-05 - -5.71534336268e-06 = 5.34336422443e-05
// Expected Z = 00111000011000000001110111110000
#10 a = 32'b00111000010010000010010100100010; b = 32'b10110110101111111100011001101101; operation = 1'b1; $display("%b", result);

// TEST #836
// -9.39211615146e-05 - 6.739357295e-05 = -0.000161314734465
// Expected Z = 10111001001010010010011010011000
#10 a = 32'b10111000110001001111011110001010; b = 32'b00111000100011010101010110100110; operation = 1'b1; $display("%b", result);

// TEST #837
// -7.42797733412e-05 - 7.38688197009e-06 = -8.16666553112e-05
// Expected Z = 10111000101010110100010001110100
#10 a = 32'b10111000100110111100011010100110; b = 32'b00110110111101111101110011010101; operation = 1'b1; $display("%b", result);

// TEST #838
// -7.25165029392e-05 - 1.31673324866e-05 = -8.56838354258e-05
// Expected Z = 10111000101100111011000100101001
#10 a = 32'b10111000100110000001010000000000; b = 32'b00110111010111001110100101000011; operation = 1'b1; $display("%b", result);

// TEST #839
// -5.12421437076e-05 - 3.29876034702e-05 = -8.42297471778e-05
// Expected Z = 10111000101100001010010010000000
#10 a = 32'b10111000010101101110110011010101; b = 32'b00111000000010100101110000101011; operation = 1'b1; $display("%b", result);

// TEST #840
// -4.38029684103e-05 + -1.42644498453e-05 = -5.80674182555e-05
// Expected Z = 10111000011100111000110101101010
#10 a = 32'b10111000001101111011100100010100; b = 32'b10110111011011110101000101011000; operation = 1'b0; $display("%b", result);

// TEST #841
// -9.47212378355e-05 + 2.49939871786e-05 = -6.97272506569e-05
// Expected Z = 10111000100100100011101010001000
#10 a = 32'b10111000110001101010010100010100; b = 32'b00110111110100011010101000101110; operation = 1'b0; $display("%b", result);

// TEST #842
// 9.352009109e-06 - -7.27180913818e-05 = 8.20701004908e-05
// Expected Z = 00111000101011000001110100001101
#10 a = 32'b00110111000111001110011010010011; b = 32'b10111000100110001000000000111010; operation = 1'b1; $display("%b", result);

// TEST #843
// 1.45595698141e-05 - 1.42243751226e-05 = 3.35194691471e-07
// Expected Z = 00110100101100111111010011001111
#10 a = 32'b00110111011101000100010011100000; b = 32'b00110111011011101010010100111010; operation = 1'b1; $display("%b", result);

// TEST #844
// -1.88362147876e-05 + 1.92232251883e-05 = 3.87010400669e-07
// Expected Z = 00110100110011111100011001001110
#10 a = 32'b10110111100111100000001001110111; b = 32'b00110111101000010100000110010000; operation = 1'b0; $display("%b", result);

// TEST #845
// 4.22440788395e-06 + 2.34956207412e-05 = 2.77200286251e-05
// Expected Z = 00110111111010001000100001001111
#10 a = 32'b00110110100011011011111101100011; b = 32'b00110111110001010001100001110110; operation = 1'b0; $display("%b", result);

// TEST #846
// -9.46341807511e-05 - -5.05743450118e-05 = -4.40598357394e-05
// Expected Z = 10111000001110001100110011100011
#10 a = 32'b10111000110001100111011001010111; b = 32'b10111000010101000001111111001010; operation = 1'b1; $display("%b", result);

// TEST #847
// 7.37575934458e-05 - 2.4968427126e-05 = 4.87891663198e-05
// Expected Z = 00111000010011001010001011111000
#10 a = 32'b00111000100110101010111001001110; b = 32'b00110111110100010111001101001010; operation = 1'b1; $display("%b", result);

// TEST #848
// 9.00115392273e-05 + -4.88397650165e-05 = 4.11717742109e-05
// Expected Z = 00111000001011001010111111011011
#10 a = 32'b00111000101111001100010010010100; b = 32'b10111000010011001101100101001100; operation = 1'b0; $display("%b", result);

// TEST #849
// 2.01175764353e-05 + 6.31199144646e-05 = 8.32374908999e-05
// Expected Z = 00111000101011101000111111001010
#10 a = 32'b00110111101010001100001000101011; b = 32'b00111000100001000101111100111111; operation = 1'b0; $display("%b", result);

// TEST #850
// -9.8150746416e-05 + 2.04951177514e-05 = -7.76556286646e-05
// Expected Z = 10111000101000101101101100001100
#10 a = 32'b10111000110011011101011001001000; b = 32'b00110111101010111110110011101110; operation = 1'b0; $display("%b", result);

// TEST #851
// 2.70233813081e-05 + 1.35827264002e-05 = 4.06061077083e-05
// Expected Z = 00111000001010100101000001111010
#10 a = 32'b00110111111000101011000001000101; b = 32'b00110111011000111110000101011110; operation = 1'b0; $display("%b", result);

// TEST #852
// 7.36040977672e-05 - -2.21447506269e-05 = 9.57488483942e-05
// Expected Z = 00111000110010001100110011000110
#10 a = 32'b00111000100110100101101111100110; b = 32'b10110111101110011100001101111101; operation = 1'b1; $display("%b", result);

// TEST #853
// 5.29378311017e-05 - -9.95893381987e-05 = 0.0001525271693
// Expected Z = 00111001000111111110111110110011
#10 a = 32'b00111000010111100000100110010000; b = 32'b10111000110100001101101010011110; operation = 1'b1; $display("%b", result);

// TEST #854
// -9.57285963707e-05 - -4.74937125949e-05 = -4.82348837758e-05
// Expected Z = 10111000010010100100111111010000
#10 a = 32'b10111000110010001100000111100110; b = 32'b10111000010001110011001111111100; operation = 1'b1; $display("%b", result);

// TEST #855
// 8.35096308671e-05 - -4.24616655792e-05 = 0.000125971296446
// Expected Z = 00111001000001000001011100101010
#10 a = 32'b00111000101011110010000111100100; b = 32'b10111000001100100001100011011110; operation = 1'b1; $display("%b", result);

// TEST #856
// -8.5333307111e-05 - 4.12968729906e-05 = -0.000126630180102
// Expected Z = 10111001000001001100100000001000
#10 a = 32'b10111000101100101111010011111000; b = 32'b00111000001011010011011000101110; operation = 1'b1; $display("%b", result);

// TEST #857
// 8.95014780074e-05 - 4.83073421785e-05 = 4.11941358288e-05
// Expected Z = 00111000001011001100011111011110
#10 a = 32'b00111000101110111011001010111101; b = 32'b00111000010010101001110110011101; operation = 1'b1; $display("%b", result);

// TEST #858
// -8.82580333703e-05 - -9.51016868135e-05 = 6.84365344321e-06
// Expected Z = 00110110111001011010001010001001
#10 a = 32'b10111000101110010001011100101100; b = 32'b10111000110001110111000101010100; operation = 1'b1; $display("%b", result);

// TEST #859
// 2.02906193921e-05 - -9.52224219364e-05 = 0.000115513041328
// Expected Z = 00111000111100100011111110011000
#10 a = 32'b00110111101010100011010111000110; b = 32'b10111000110001111011001000100110; operation = 1'b1; $display("%b", result);

// TEST #860
// -2.16214093708e-05 + 7.78972261015e-05 = 5.62758167306e-05
// Expected Z = 00111000011011000000100110110011
#10 a = 32'b10110111101101010101111110100000; b = 32'b00111000101000110101110011000001; operation = 1'b0; $display("%b", result);

// TEST #861
// 7.2613070054e-05 + 2.89724622598e-05 = 0.000101585532314
// Expected Z = 00111000110101010000101001010001
#10 a = 32'b00111000100110000100011111011000; b = 32'b00110111111100110000100111100100; operation = 1'b0; $display("%b", result);

// TEST #862
// -7.63674428907e-05 - 1.07678663045e-06 = -7.74442295211e-05
// Expected Z = 10111000101000100110100110001110
#10 a = 32'b10111000101000000010011101110101; b = 32'b00110101100100001000011000011011; operation = 1'b1; $display("%b", result);

// TEST #863
// 1.26005019984e-05 + 8.73235944664e-05 = 9.99240964648e-05
// Expected Z = 00111000110100011000111001010111
#10 a = 32'b00110111010100110110011010111110; b = 32'b00111000101101110010000101111111; operation = 1'b0; $display("%b", result);

// TEST #864
// -4.2370719096e-05 - 2.61942868723e-05 = -6.85650059684e-05
// Expected Z = 10111000100011111100101010001111
#10 a = 32'b10111000001100011011011100110111; b = 32'b00110111110110111011101111001101; operation = 1'b1; $display("%b", result);

// TEST #865
// -3.14794434326e-05 - 5.60369119679e-05 = -8.75163554005e-05
// Expected Z = 10111000101101111000100011111100
#10 a = 32'b10111000000001000000100011001100; b = 32'b00111000011010110000100100101101; operation = 1'b1; $display("%b", result);

// TEST #866
// -4.9440900057e-05 - -6.1406232494e-05 = 1.1965332437e-05
// Expected Z = 00110111010010001011111010110110
#10 a = 32'b10111000010011110101111011000011; b = 32'b10111000100000001100011100111000; operation = 1'b1; $display("%b", result);

// TEST #867
// -2.49592517909e-05 + 1.48684036936e-06 = -2.34724114215e-05
// Expected Z = 10110111110001001110011010011111
#10 a = 32'b10110111110100010101111110010110; b = 32'b00110101110001111000111101110010; operation = 1'b0; $display("%b", result);

// TEST #868
// 8.87702579203e-05 + -1.40541144947e-05 = 7.47161434256e-05
// Expected Z = 00111000100111001011000011101101
#10 a = 32'b00111000101110100010101000101011; b = 32'b10110111011010111100100111110110; operation = 1'b0; $display("%b", result);

// TEST #869
// -9.32065171979e-05 - -6.79890190793e-06 = -8.640761529e-05
// Expected Z = 10111000101101010011010110111100
#10 a = 32'b10111000110000110111011111011110; b = 32'b10110110111001000010001000011111; operation = 1'b1; $display("%b", result);

// TEST #870
// 6.76746886476e-05 - -3.75591784575e-05 = 0.000105233867105
// Expected Z = 00111000110111001011000100000001
#10 a = 32'b00111000100011011110110010010010; b = 32'b10111000000111011000100011011100; operation = 1'b1; $display("%b", result);

// TEST #871
// 2.17276054076e-05 - 1.10263576803e-05 = 1.07012477273e-05
// Expected Z = 00110111001100111000100110000010
#10 a = 32'b00110111101101100100001110101101; b = 32'b00110111001110001111110111011000; operation = 1'b1; $display("%b", result);

// TEST #872
// 6.51498175605e-05 - 3.74496538735e-05 = 2.7700163687e-05
// Expected Z = 00110111111010000101110110100110
#10 a = 32'b00111000100010001010000100001011; b = 32'b00111000000111010001001101000010; operation = 1'b1; $display("%b", result);

// TEST #873
// -3.45075530553e-05 - 8.56481433112e-05 = -0.000120155696366
// Expected Z = 10111000111110111111110000011001
#10 a = 32'b10111000000100001011110000110100; b = 32'b00111000101100111001110111111111; operation = 1'b1; $display("%b", result);

// TEST #874
// 7.00154174448e-06 + -6.74093256878e-05 = -6.04077839433e-05
// Expected Z = 10111000011111010101111001011101
#10 a = 32'b00110110111010101110111011001001; b = 32'b10111000100011010101111000011011; operation = 1'b0; $display("%b", result);

// TEST #875
// -4.25686702618e-05 - -4.17050233208e-05 = -8.63646941008e-07
// Expected Z = 10110101011001111101010101011110
#10 a = 32'b10111000001100101000101111000011; b = 32'b10111000001011101110110001101110; operation = 1'b1; $display("%b", result);

// TEST #876
// 4.87913038357e-05 + 4.68333503719e-05 = 9.56246542075e-05
// Expected Z = 00111000110010001000101000011000
#10 a = 32'b00111000010011001010010101000011; b = 32'b00111000010001000110111011101101; operation = 1'b0; $display("%b", result);

// TEST #877
// -1.24202100027e-07 + -3.29995213298e-05 = -3.31237234298e-05
// Expected Z = 10111000000010101110111001010100
#10 a = 32'b10110100000001010101110001101010; b = 32'b10111000000010100110100011110111; operation = 1'b0; $display("%b", result);

// TEST #878
// -6.50044886093e-05 - -3.69565369332e-05 = -2.80479516761e-05
// Expected Z = 10110111111010110100100010000101
#10 a = 32'b10111000100010000101001100000101; b = 32'b10111000000110110000000111001000; operation = 1'b1; $display("%b", result);

// TEST #879
// 5.35958028993e-05 + -3.7464698518e-05 = 1.61311043813e-05
// Expected Z = 00110111100001110101000101001000
#10 a = 32'b00111000011000001100110000001110; b = 32'b10111000000111010010001101101010; operation = 1'b0; $display("%b", result);

// TEST #880
// 6.79193790151e-05 - 4.42555955305e-05 = 2.36637834846e-05
// Expected Z = 00110111110001101000000110010111
#10 a = 32'b00111000100011100110111111110000; b = 32'b00111000001110011001111100010101; operation = 1'b1; $display("%b", result);

// TEST #881
// -9.85161016894e-05 - -9.18469450154e-05 = -6.66915667396e-06
// Expected Z = 10110110110111111100011110011111
#10 a = 32'b10111000110011101001101001101110; b = 32'b10111000110000001001110111110100; operation = 1'b1; $display("%b", result);

// TEST #882
// -1.05123478161e-05 - -8.76376719993e-07 = -9.63597109606e-06
// Expected Z = 10110111001000011010101000101110
#10 a = 32'b10110111001100000101111000110001; b = 32'b10110101011010110100000000100110; operation = 1'b1; $display("%b", result);

// TEST #883
// 5.47484423864e-05 + 2.99162446854e-05 = 8.46646870718e-05
// Expected Z = 00111000101100011000111000000010
#10 a = 32'b00111000011001011010000110110001; b = 32'b00110111111110101111010010100101; operation = 1'b0; $display("%b", result);

// TEST #884
// 7.86559820543e-05 - 2.62464119259e-05 = 5.24095701284e-05
// Expected Z = 00111000010110111101001001011001
#10 a = 32'b00111000101001001111010000011100; b = 32'b00110111110111000010101110111110; operation = 1'b1; $display("%b", result);

// TEST #885
// -7.38355428399e-06 + 6.47088539302e-05 = 5.73252996462e-05
// Expected Z = 00111000011100000111000010010010
#10 a = 32'b10110110111101111100000001000000; b = 32'b00111000100001111011010001001101; operation = 1'b0; $display("%b", result);

// TEST #886
// 9.79161159333e-06 + -6.23817866854e-05 = -5.25901750921e-05
// Expected Z = 10111000010111001001010001000101
#10 a = 32'b00110111001001000100011010100111; b = 32'b10111000100000101101001011110111; operation = 1'b0; $display("%b", result);

// TEST #887
// -2.9308092131e-05 - -5.74460234316e-05 = 2.81379313007e-05
// Expected Z = 00110111111011000000100110111111
#10 a = 32'b10110111111101011101101010100110; b = 32'b10111000011100001111001000110011; operation = 1'b1; $display("%b", result);

// TEST #888
// 5.74089929291e-05 - -2.70043752336e-05 = 8.44133681627e-05
// Expected Z = 00111000101100010000011100010101
#10 a = 32'b00111000011100001100101001110000; b = 32'b10110111111000101000011101110100; operation = 1'b1; $display("%b", result);

// TEST #889
// -9.97449070569e-05 - -4.10499055671e-05 = -5.86950014898e-05
// Expected Z = 10111000011101100010111101000111
#10 a = 32'b10111000110100010010111000100100; b = 32'b10111000001011000010110100000000; operation = 1'b1; $display("%b", result);

// TEST #890
// -7.80159634247e-05 + 7.92093694605e-05 = 1.19340603575e-06
// Expected Z = 00110101101000000010110100011111
#10 a = 32'b10111000101000111001110010000000; b = 32'b00111000101001100001110100110101; operation = 1'b0; $display("%b", result);

// TEST #891
// -1.77274053889e-05 + -2.5206947778e-05 = -4.29343531669e-05
// Expected Z = 10111000001101000001010001101001
#10 a = 32'b10110111100101001011010101010000; b = 32'b10110111110100110111001110000010; operation = 1'b0; $display("%b", result);

// TEST #892
// 6.46923966326e-05 + -6.92448495974e-05 = -4.55245296481e-06
// Expected Z = 10110110100110001100000101000110
#10 a = 32'b00111000100001111010101101110111; b = 32'b10111000100100010011011110001100; operation = 1'b0; $display("%b", result);

// TEST #893
// 3.53959083632e-05 - 4.41908242338e-05 = -8.79491587056e-06
// Expected Z = 10110111000100111000110111100000
#10 a = 32'b00111000000101000111011000010001; b = 32'b00111000001110010101100110001001; operation = 1'b1; $display("%b", result);

// TEST #894
// 3.83124900751e-05 + 7.80503954226e-05 = 0.000116362885498
// Expected Z = 00111000111101000000011111011001
#10 a = 32'b00111000001000001011000110111001; b = 32'b00111000101000111010111011111101; operation = 1'b0; $display("%b", result);

// TEST #895
// 3.65511547245e-05 - -4.58578645661e-05 = 8.24090192906e-05
// Expected Z = 00111000101011001101001100000001
#10 a = 32'b00111000000110010100111010000001; b = 32'b10111000010000000101011110000010; operation = 1'b1; $display("%b", result);

// TEST #896
// -9.80624515271e-05 + -3.86326094773e-05 = -0.000136695061004
// Expected Z = 10111001000011110101010111001101
#10 a = 32'b10111000110011011010011011100001; b = 32'b10111000001000100000100101110011; operation = 1'b0; $display("%b", result);

// TEST #897
// -3.80734190187e-05 + -7.86485973054e-06 = -4.59382787492e-05
// Expected Z = 10111000010000001010110111011010
#10 a = 32'b10111000000111111011000100000110; b = 32'b10110111000000111111001101010001; operation = 1'b0; $display("%b", result);

// TEST #898
// 6.44706802045e-05 - -3.33659755399e-05 = 9.78366557444e-05
// Expected Z = 00111000110011010010110110101000
#10 a = 32'b00111000100001110011010001101111; b = 32'b10111000000010111111001001110010; operation = 1'b1; $display("%b", result);

// TEST #899
// -8.03812348923e-05 + -7.21284398497e-05 = -0.000152509674742
// Expected Z = 10111001000111111110101100000001
#10 a = 32'b10111000101010001001001001011001; b = 32'b10111000100101110100001110101001; operation = 1'b0; $display("%b", result);

// TEST #900
// -4.36997421696e-05 - -3.05073137461e-05 = -1.31924284235e-05
// Expected Z = 10110111010111010101010100001100
#10 a = 32'b10111000001101110100101000111110; b = 32'b10110111111111111110100111110101; operation = 1'b1; $display("%b", result);

// TEST #901
// -229574.197877 - 84360.0403897 = -313934.238267
// Expected Z = 11001000100110010100100111001000
#10 a = 32'b11001000011000000011000110001101; b = 32'b01000111101001001100010000000101; operation = 1'b1; $display("%b", result);

// TEST #902
// -373766.567662 - 158750.547368 = -532517.11503
// Expected Z = 11001001000000100000001001010010
#10 a = 32'b11001000101101101000000011010010; b = 32'b01001000000110110000011110100011; operation = 1'b1; $display("%b", result);

// TEST #903
// -884246.672281 + -25396.2852957 = -909642.957577
// Expected Z = 11001001010111100001010010101111
#10 a = 32'b11001001010101111110000101101011; b = 32'b11000110110001100110100010010010; operation = 1'b0; $display("%b", result);

// TEST #904
// -571742.678139 - -313182.175186 = -258560.502954
// Expected Z = 11001000011111001000000000100000
#10 a = 32'b11001001000010111001010111101011; b = 32'b11001000100110001110101111000110; operation = 1'b1; $display("%b", result);

// TEST #905
// -676152.853814 + -519215.809897 = -1195368.66371
// Expected Z = 11001001100100011110101101000101
#10 a = 32'b11001001001001010001001110001110; b = 32'b11001000111111011000010111111010; operation = 1'b0; $display("%b", result);

// TEST #906
// 699821.938929 - 193087.505903 = 506734.433026
// Expected Z = 01001000111101110110110111001110
#10 a = 32'b01001001001010101101101011011111; b = 32'b01001000001111001000111111100000; operation = 1'b1; $display("%b", result);

// TEST #907
// 336903.338014 + 72147.6618781 = 409050.999892
// Expected Z = 01001000110001111011101101100000
#10 a = 32'b01001000101001001000000011101011; b = 32'b01000111100011001110100111010101; operation = 1'b0; $display("%b", result);

// TEST #908
// 697219.56897 - -896872.625164 = 1594092.19413
// Expected Z = 01001001110000101001011101100010
#10 a = 32'b01001001001010100011100000111001; b = 32'b11001001010110101111011010001010; operation = 1'b1; $display("%b", result);

// TEST #909
// -891730.228887 - 712858.694148 = -1604588.92303
// Expected Z = 11001001110000111101111101100111
#10 a = 32'b11001001010110011011010100100100; b = 32'b01001001001011100000100110101011; operation = 1'b1; $display("%b", result);

// TEST #910
// 226236.392918 + -31558.6740998 = 194677.718819
// Expected Z = 01001000001111100001110101101110
#10 a = 32'b01001000010111001110111100011001; b = 32'b11000110111101101000110101011001; operation = 1'b0; $display("%b", result);

// TEST #911
// -311807.411871 - -941879.515736 = 630072.103865
// Expected Z = 01001001000110011101001110000010
#10 a = 32'b11001000100110000011111111101101; b = 32'b11001001011001011111001101111000; operation = 1'b1; $display("%b", result);

// TEST #912
// -258900.653621 + -878184.261404 = -1137084.91503
// Expected Z = 11001001100010101100110111100111
#10 a = 32'b11001000011111001101010100101010; b = 32'b11001001010101100110011010000100; operation = 1'b0; $display("%b", result);

// TEST #913
// 436101.907666 - 534243.952631 = -98142.0449654
// Expected Z = 11000111101111111010111100000110
#10 a = 32'b01001000110101001111000010111101; b = 32'b01001001000000100110111000111111; operation = 1'b1; $display("%b", result);

// TEST #914
// 153820.494071 - 614212.262382 = -460391.768311
// Expected Z = 11001000111000001100110011111001
#10 a = 32'b01001000000101100011011100100000; b = 32'b01001001000101011111010001000100; operation = 1'b1; $display("%b", result);

// TEST #915
// 404284.373674 - 242036.271929 = 162248.101746
// Expected Z = 01001000000111100111001000000111
#10 a = 32'b01001000110001010110011110001100; b = 32'b01001000011011000101110100010001; operation = 1'b1; $display("%b", result);

// TEST #916
// 727423.196638 + 876909.744588 = 1604332.94123
// Expected Z = 01001001110000111101011101101000
#10 a = 32'b01001001001100011001011111110011; b = 32'b01001001010101100001011011011100; operation = 1'b0; $display("%b", result);

// TEST #917
// -421731.514826 + -965612.915196 = -1387344.43002
// Expected Z = 11001001101010010101101010000011
#10 a = 32'b11001000110011011110110001110000; b = 32'b11001001011010111011111011001111; operation = 1'b0; $display("%b", result);

// TEST #918
// 104559.377958 + -792244.742373 = -687685.364415
// Expected Z = 11001001001001111110010001010110
#10 a = 32'b01000111110011000011011110110000; b = 32'b11001001010000010110101101001100; operation = 1'b0; $display("%b", result);

// TEST #919
// -630415.247559 + -481920.228751 = -1112335.47631
// Expected Z = 11001001100001111100100001111100
#10 a = 32'b11001001000110011110100011110100; b = 32'b11001000111010110101000000000111; operation = 1'b0; $display("%b", result);

// TEST #920
// -618111.251678 + 756056.972746 = 137945.721068
// Expected Z = 01001000000001101011011001101110
#10 a = 32'b11001001000101101110011111110100; b = 32'b01001001001110001001010110010000; operation = 1'b0; $display("%b", result);

// TEST #921
// 446106.887599 + -833512.46124 = -387405.573641
// Expected Z = 11001000101111010010100110110010
#10 a = 32'b01001000110110011101001101011100; b = 32'b11001001010010110111111010000111; operation = 1'b0; $display("%b", result);

// TEST #922
// -495445.631984 + -868851.688365 = -1364297.32035
// Expected Z = 11001001101001101000101001001011
#10 a = 32'b11001000111100011110101010110100; b = 32'b11001001010101000001111100111011; operation = 1'b0; $display("%b", result);

// TEST #923
// 91323.2418801 + -409621.067091 = -318297.825211
// Expected Z = 11001000100110110110101100111010
#10 a = 32'b01000111101100100101110110011111; b = 32'b11001000110010000000001010100010; operation = 1'b0; $display("%b", result);

// TEST #924
// 738184.326099 + -670707.002984 = 67477.3231149
// Expected Z = 01000111100000111100101010101001
#10 a = 32'b01001001001101000011100010000101; b = 32'b11001001001000111011111100110000; operation = 1'b0; $display("%b", result);

// TEST #925
// 242170.46398 + -876209.026315 = -634038.562335
// Expected Z = 11001001000110101100101101101001
#10 a = 32'b01001000011011000111111010011110; b = 32'b11001001010101011110101100010000; operation = 1'b0; $display("%b", result);

// TEST #926
// -724134.726635 + 862949.846079 = 138815.119444
// Expected Z = 01001000000001111000111111001000
#10 a = 32'b11001001001100001100101001101100; b = 32'b01001001010100101010111001011110; operation = 1'b0; $display("%b", result);

// TEST #927
// 561181.34343 - 120991.621969 = 440189.721461
// Expected Z = 01001000110101101110111110110111
#10 a = 32'b01001001000010010000000111010101; b = 32'b01000111111011000100111111010000; operation = 1'b1; $display("%b", result);

// TEST #928
// -730813.01544 - -438244.971829 = -292568.04361
// Expected Z = 11001000100011101101101100000001
#10 a = 32'b11001001001100100110101111010000; b = 32'b11001000110101011111110010011111; operation = 1'b1; $display("%b", result);

// TEST #929
// -12160.3463607 + -465093.212667 = -477253.559028
// Expected Z = 11001000111010010000100010110010
#10 a = 32'b11000110001111100000000101100011; b = 32'b11001000111000110001100010100111; operation = 1'b0; $display("%b", result);

// TEST #930
// -114165.463989 - 853696.913874 = -967862.377863
// Expected Z = 11001001011011000100101101100110
#10 a = 32'b11000111110111101111101010111011; b = 32'b01001001010100000110110000001111; operation = 1'b1; $display("%b", result);

// TEST #931
// 896133.825831 + -745767.16476 = 150366.661071
// Expected Z = 01001000000100101101011110101010
#10 a = 32'b01001001010110101100100001011101; b = 32'b11001001001101100001001001110011; operation = 1'b0; $display("%b", result);

// TEST #932
// 623606.921408 + 613344.737066 = 1236951.65847
// Expected Z = 01001001100101101111111010111101
#10 a = 32'b01001001000110000011111101101111; b = 32'b01001001000101011011111000001100; operation = 1'b0; $display("%b", result);

// TEST #933
// 382551.003613 + 316758.796343 = 699309.799956
// Expected Z = 01001001001010101011101011011101
#10 a = 32'b01001000101110101100101011100000; b = 32'b01001000100110101010101011011001; operation = 1'b0; $display("%b", result);

// TEST #934
// 88417.1309438 + 64166.605305 = 152583.736249
// Expected Z = 01001000000101010000000111101111
#10 a = 32'b01000111101011001011000010010001; b = 32'b01000111011110101010011010011011; operation = 1'b0; $display("%b", result);

// TEST #935
// -220484.69853 + -476558.957512 = -697043.656042
// Expected Z = 11001001001010100010110100111010
#10 a = 32'b11001000010101110101000100101101; b = 32'b11001000111010001011000111011111; operation = 1'b0; $display("%b", result);

// TEST #936
// 636619.566206 + 438804.356963 = 1075423.92317
// Expected Z = 01001001100000110100011011111111
#10 a = 32'b01001001000110110110110010111001; b = 32'b01001000110101100100001010001011; operation = 1'b0; $display("%b", result);

// TEST #937
// 867924.265591 - 606224.877085 = 261699.388507
// Expected Z = 01001000011111111001000011011001
#10 a = 32'b01001001010100111110010101000100; b = 32'b01001001000101000000000100001110; operation = 1'b1; $display("%b", result);

// TEST #938
// -212867.43009 + -156704.190847 = -369571.620937
// Expected Z = 11001000101101000111010001110100
#10 a = 32'b11001000010011111110000011011100; b = 32'b11001000000110010000100000001100; operation = 1'b0; $display("%b", result);

// TEST #939
// 339173.452045 - 652324.042409 = -313150.590364
// Expected Z = 11001000100110001110011111010011
#10 a = 32'b01001000101001011001110010101110; b = 32'b01001001000111110100001001000001; operation = 1'b1; $display("%b", result);

// TEST #940
// 674194.016899 - -44108.9130851 = 718302.929984
// Expected Z = 01001001001011110101110111101111
#10 a = 32'b01001001001001001001100100100000; b = 32'b11000111001011000100110011101010; operation = 1'b1; $display("%b", result);

// TEST #941
// -900956.391554 - -894096.243827 = -6860.14772658
// Expected Z = 11000101110101100110000100101111
#10 a = 32'b11001001010110111111010111000110; b = 32'b11001001010110100100100100000100; operation = 1'b1; $display("%b", result);

// TEST #942
// 218748.741317 - -69729.8537217 = 288478.595039
// Expected Z = 01001000100011001101101111010011
#10 a = 32'b01001000010101011001111100101111; b = 32'b11000111100010000011000011101101; operation = 1'b1; $display("%b", result);

// TEST #943
// -954632.927732 - 412997.025951 = -1367629.95368
// Expected Z = 11001001101001101111001001110000
#10 a = 32'b11001001011010010001000010001111; b = 32'b01001000110010011010100010100001; operation = 1'b1; $display("%b", result);

// TEST #944
// -107050.01544 - -458160.715713 = 351110.700274
// Expected Z = 01001000101010110111000011010110
#10 a = 32'b11000111110100010001010100000010; b = 32'b11001000110111111011011000010111; operation = 1'b1; $display("%b", result);

// TEST #945
// -940061.648305 + -17314.6994821 = -957376.347787
// Expected Z = 11001001011010011011110000000110
#10 a = 32'b11001001011001011000000111011010; b = 32'b11000110100001110100010101100110; operation = 1'b0; $display("%b", result);

// TEST #946
// 488647.039104 - -377916.286205 = 866563.325308
// Expected Z = 01001001010100111001000000110101
#10 a = 32'b01001000111011101001100011100001; b = 32'b11001000101110001000011110001001; operation = 1'b1; $display("%b", result);

// TEST #947
// 508428.375999 - 354078.854406 = 154349.521593
// Expected Z = 01001000000101101011101101100001
#10 a = 32'b01001000111110000100000110001100; b = 32'b01001000101011001110001111011011; operation = 1'b1; $display("%b", result);

// TEST #948
// -346304.080417 - 304623.35042 = -650927.430837
// Expected Z = 11001001000111101110101011110111
#10 a = 32'b11001000101010010001100000000011; b = 32'b01001000100101001011110111101011; operation = 1'b1; $display("%b", result);

// TEST #949
// 980358.092967 - -922464.409792 = 1902822.50276
// Expected Z = 01001001111010000100011100110100
#10 a = 32'b01001001011011110101100001100001; b = 32'b11001001011000010011011000000111; operation = 1'b1; $display("%b", result);

// TEST #950
// -398419.647724 - -337805.465397 = -60614.1823278
// Expected Z = 11000111011011001100011000101111
#10 a = 32'b11001000110000101000101001110101; b = 32'b11001000101001001111000110101111; operation = 1'b1; $display("%b", result);

// TEST #951
// -934976.561438 - 19930.5976858 = -954907.159124
// Expected Z = 11001001011010010010000110110011
#10 a = 32'b11001001011001000100010000001001; b = 32'b01000110100110111011010100110010; operation = 1'b1; $display("%b", result);

// TEST #952
// -184769.843686 + 176522.032937 = -8247.81074989
// Expected Z = 11000110000000001101111100111110
#10 a = 32'b11001000001101000111000001110110; b = 32'b01001000001011000110001010000010; operation = 1'b0; $display("%b", result);

// TEST #953
// -387993.860543 - 188678.892578 = -576672.753121
// Expected Z = 11001001000011001100101000001100
#10 a = 32'b11001000101111010111001100111100; b = 32'b01001000001110000100000110111001; operation = 1'b1; $display("%b", result);

// TEST #954
// -635338.007592 + -596526.660535 = -1231864.66813
// Expected Z = 11001001100101100101111111000101
#10 a = 32'b11001001000110110001110010100000; b = 32'b11001001000100011010001011101011; operation = 1'b0; $display("%b", result);

// TEST #955
// 210634.218301 + 880346.177197 = 1090980.3955
// Expected Z = 01001001100001010010110100100011
#10 a = 32'b01001000010011011011001010001110; b = 32'b01001001010101101110110110100011; operation = 1'b0; $display("%b", result);

// TEST #956
// -920441.762717 - -223760.614229 = -696681.148488
// Expected Z = 11001001001010100001011010010010
#10 a = 32'b11001001011000001011011110011100; b = 32'b11001000010110101000010000100111; operation = 1'b1; $display("%b", result);

// TEST #957
// -701502.069369 + -553854.314024 = -1255356.38339
// Expected Z = 11001001100110010011110111100011
#10 a = 32'b11001001001010110100001111100001; b = 32'b11001001000001110011011111100101; operation = 1'b0; $display("%b", result);

// TEST #958
// 397294.005294 + 397448.043865 = 794742.049159
// Expected Z = 01001001010000100000011101100001
#10 a = 32'b01001000110000011111110111000000; b = 32'b01001000110000100001000100000001; operation = 1'b0; $display("%b", result);

// TEST #959
// 553741.016234 + -379058.772113 = 174682.244121
// Expected Z = 01001000001010101001011010010000
#10 a = 32'b01001001000001110011000011010000; b = 32'b11001000101110010001011001011001; operation = 1'b0; $display("%b", result);

// TEST #960
// 459196.198378 - -941455.209795 = 1400651.40817
// Expected Z = 01001001101010101111101001011011
#10 a = 32'b01001000111000000011011110000110; b = 32'b11001001011001011101100011110011; operation = 1'b1; $display("%b", result);

// TEST #961
// 209747.183118 + -781774.192018 = -572027.0089
// Expected Z = 11001001000010111010011110110000
#10 a = 32'b01001000010011001101010011001100; b = 32'b11001001001111101101110011100011; operation = 1'b0; $display("%b", result);

// TEST #962
// 420507.014275 + 617574.788526 = 1038081.8028
// Expected Z = 01001001011111010111000000011101
#10 a = 32'b01001000110011010101001101100000; b = 32'b01001001000101101100011001101101; operation = 1'b0; $display("%b", result);

// TEST #963
// 302872.442795 - -229526.643478 = 532399.086273
// Expected Z = 01001001000000011111101011110001
#10 a = 32'b01001000100100111110001100001110; b = 32'b11001000011000000010010110101001; operation = 1'b1; $display("%b", result);

// TEST #964
// 314358.716133 - 671862.595611 = -357503.879478
// Expected Z = 11001000101011101000111111111100
#10 a = 32'b01001000100110010111111011010111; b = 32'b01001001001001000000011101101010; operation = 1'b1; $display("%b", result);

// TEST #965
// -702829.186543 + -963049.204893 = -1665878.39144
// Expected Z = 11001001110010110101101010110011
#10 a = 32'b11001001001010111001011011010011; b = 32'b11001001011010110001111010010011; operation = 1'b0; $display("%b", result);

// TEST #966
// -976211.646702 + -963831.673123 = -1940043.31982
// Expected Z = 11001001111011001101001001011011
#10 a = 32'b11001001011011100101010100111010; b = 32'b11001001011010110100111101111011; operation = 1'b0; $display("%b", result);

// TEST #967
// -160716.408691 - 666097.083968 = -826813.492659
// Expected Z = 11001001010010011101101111011000
#10 a = 32'b11001000000111001111001100011010; b = 32'b01001001001000101001111100010001; operation = 1'b1; $display("%b", result);

// TEST #968
// 785347.480403 - 438043.037678 = 347304.442725
// Expected Z = 01001000101010011001010100001110
#10 a = 32'b01001001001111111011110000111000; b = 32'b01001000110101011110001101100001; operation = 1'b1; $display("%b", result);

// TEST #969
// -718645.839863 + 46479.5042995 = -672166.335564
// Expected Z = 11001001001001000001101001100101
#10 a = 32'b11001001001011110111001101011101; b = 32'b01000111001101011000111110000001; operation = 1'b0; $display("%b", result);

// TEST #970
// -468684.835005 + 834543.54486 = 365858.709855
// Expected Z = 01001000101100101010010001010111
#10 a = 32'b11001000111001001101100110011011; b = 32'b01001001010010111011111011111001; operation = 1'b0; $display("%b", result);

// TEST #971
// 495817.11646 + -906369.544238 = -410552.427778
// Expected Z = 11001000110010000111011100001110
#10 a = 32'b01001000111100100001100100100100; b = 32'b11001001010111010100100000011001; operation = 1'b0; $display("%b", result);

// TEST #972
// -810671.259803 - 662620.16145 = -1473291.42125
// Expected Z = 11001001101100111101100001011011
#10 a = 32'b11001001010001011110101011110100; b = 32'b01001001001000011100010111000011; operation = 1'b1; $display("%b", result);

// TEST #973
// 979476.684126 + 30926.4472771 = 1010403.1314
// Expected Z = 01001001011101101010111000110010
#10 a = 32'b01001001011011110010000101001011; b = 32'b01000110111100011001110011100101; operation = 1'b0; $display("%b", result);

// TEST #974
// 225577.992997 + 794.984148208 = 226372.977145
// Expected Z = 01001000010111010001000100111111
#10 a = 32'b01001000010111000100101010000000; b = 32'b01000100010001101011111011111100; operation = 1'b0; $display("%b", result);

// TEST #975
// 321962.665843 + -599970.920715 = -278008.254872
// Expected Z = 11001000100001111011111100001000
#10 a = 32'b01001000100111010011010101010101; b = 32'b11001001000100100111101000101111; operation = 1'b0; $display("%b", result);

// TEST #976
// -297261.483741 + -25455.0224666 = -322716.506208
// Expected Z = 11001000100111011001001110010000
#10 a = 32'b11001000100100010010010110101111; b = 32'b11000110110001101101111000001100; operation = 1'b0; $display("%b", result);

// TEST #977
// -443678.728654 + 764857.737391 = 321179.008737
// Expected Z = 01001000100111001101001101100000
#10 a = 32'b11001000110110001010001111010111; b = 32'b01001001001110101011101110011100; operation = 1'b0; $display("%b", result);

// TEST #978
// -350382.008791 + 605224.112721 = 254842.10393
// Expected Z = 01001000011110001101111010000111
#10 a = 32'b11001000101010110001010111000000; b = 32'b01001001000100111100001010000010; operation = 1'b0; $display("%b", result);

// TEST #979
// -154541.511939 - 343902.141962 = -498443.653901
// Expected Z = 11001000111100110110000101110101
#10 a = 32'b11001000000101101110101101100001; b = 32'b01001000101001111110101111000101; operation = 1'b1; $display("%b", result);

// TEST #980
// -476325.2431 + 995216.878922 = 518891.635823
// Expected Z = 01001000111111010101110101110100
#10 a = 32'b11001000111010001001010010101000; b = 32'b01001001011100101111100100001110; operation = 1'b0; $display("%b", result);

// TEST #981
// -129513.548706 + -686687.801777 = -816201.350483
// Expected Z = 11001001010001110100010010010110
#10 a = 32'b11000111111111001111010011000110; b = 32'b11001001001001111010010111111101; operation = 1'b0; $display("%b", result);

// TEST #982
// -638766.995305 - 375573.322114 = -1014340.31742
// Expected Z = 11001001011101111010010001000101
#10 a = 32'b11001001000110111111001011110000; b = 32'b01001000101101110110001010101010; operation = 1'b1; $display("%b", result);

// TEST #983
// 303024.469509 - 603852.882339 = -300828.41283
// Expected Z = 11001000100100101110001110001101
#10 a = 32'b01001000100100111111011000001111; b = 32'b01001001000100110110110011001110; operation = 1'b1; $display("%b", result);

// TEST #984
// 846457.791739 - -201239.119923 = 1047696.91166
// Expected Z = 01001001011111111100100100001111
#10 a = 32'b01001001010011101010011110011101; b = 32'b11001000010001001000010111001000; operation = 1'b1; $display("%b", result);

// TEST #985
// -258476.448799 - -612776.063025 = 354299.614227
// Expected Z = 01001000101011001111111101110100
#10 a = 32'b11001000011111000110101100011101; b = 32'b11001001000101011001101010000001; operation = 1'b1; $display("%b", result);

// TEST #986
// 499385.841087 + 798167.49202 = 1297553.33311
// Expected Z = 01001001100111100110010010001011
#10 a = 32'b01001000111100111101011100111011; b = 32'b01001001010000101101110101111000; operation = 1'b0; $display("%b", result);

// TEST #987
// -752250.330106 + 562928.238547 = -189322.091558
// Expected Z = 11001000001110001110001010000110
#10 a = 32'b11001001001101111010011110100101; b = 32'b01001001000010010110111100000100; operation = 1'b0; $display("%b", result);

// TEST #988
// -838373.713041 + 666969.835642 = -171403.877398
// Expected Z = 11001000001001110110001011111000
#10 a = 32'b11001001010011001010111001011011; b = 32'b01001001001000101101010110011101; operation = 1'b0; $display("%b", result);

// TEST #989
// -649035.555146 + 99854.7491813 = -549180.805965
// Expected Z = 11001001000001100001001111001101
#10 a = 32'b11001001000111100111010010111001; b = 32'b01000111110000110000011101100000; operation = 1'b0; $display("%b", result);

// TEST #990
// 890793.174275 + -391668.67265 = 499124.501625
// Expected Z = 01001000111100111011011010010000
#10 a = 32'b01001001010110010111101010010011; b = 32'b11001000101111110011111010010110; operation = 1'b0; $display("%b", result);

// TEST #991
// 632839.150882 + 237697.167388 = 870536.31827
// Expected Z = 01001001010101001000100010000101
#10 a = 32'b01001001000110101000000001110010; b = 32'b01001000011010000010000001001011; operation = 1'b0; $display("%b", result);

// TEST #992
// -91923.4562591 - 535781.392207 = -627704.848466
// Expected Z = 11001001000110010011111110001110
#10 a = 32'b11000111101100111000100110111010; b = 32'b01001001000000101100111001010110; operation = 1'b1; $display("%b", result);

// TEST #993
// -91310.2956819 + 783271.449284 = 691961.153602
// Expected Z = 01001001001010001110111110010010
#10 a = 32'b11000111101100100101011100100110; b = 32'b01001001001111110011101001110111; operation = 1'b0; $display("%b", result);

// TEST #994
// 608537.910033 + 673797.697833 = 1282335.60787
// Expected Z = 01001001100111001000100011111101
#10 a = 32'b01001001000101001001000110011111; b = 32'b01001001001001001000000001011011; operation = 1'b0; $display("%b", result);

// TEST #995
// -139934.221644 - 446668.045732 = -586602.267377
// Expected Z = 11001001000011110011011010100100
#10 a = 32'b11001000000010001010011110001110; b = 32'b01001000110110100001100110000001; operation = 1'b1; $display("%b", result);

// TEST #996
// 735344.781899 - -511889.672085 = 1247234.45398
// Expected Z = 01001001100110000100000000010100
#10 a = 32'b01001001001100111000011100001101; b = 32'b11001000111110011111001000110110; operation = 1'b1; $display("%b", result);

// TEST #997
// -50510.0155132 + 894663.569095 = 844153.553582
// Expected Z = 01001001010011100001011110011001
#10 a = 32'b11000111010001010100111000000100; b = 32'b01001001010110100110110001111001; operation = 1'b0; $display("%b", result);

// TEST #998
// -931073.045058 - -469676.254136 = -461396.790922
// Expected Z = 11001000111000010100101010011001
#10 a = 32'b11001001011000110101000000010001; b = 32'b11001000111001010101010110001000; operation = 1'b1; $display("%b", result);

// TEST #999
// 359203.652135 + 461983.159082 = 821186.811218
// Expected Z = 01001001010010000111110000101101
#10 a = 32'b01001000101011110110010001110101; b = 32'b01001000111000011001001111100101; operation = 1'b0; $display("%b", result);

// TEST #1000
// 287625.936055 - -872985.908317 = 1160611.84437
// Expected Z = 01001001100011011010110100011111
#10 a = 32'b01001000100011000111000100111110; b = 32'b11001001010101010010000110011111; operation = 1'b1; $display("%b", result);

for(i=0; i<=10; i=i+1) begin
	#10 $display("%b", result); 
end 

#100 

#10 $finish; 

	end
      
endmodule

