`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// Create Date:    08:40:21 09/19/2012 
// Module Name:    FPMult
// Project Name: 	 Floating Point Project
// Author:			 Fredrik Brosser
//
//////////////////////////////////////////////////////////////////////////////////

module FPMult(
		A,
		B,
		Ctrl,
		P
    );
	
	// Input Ports
	input [31:0] A;
	input [31:0] B;
	input [2:0] Ctrl;
	
	// Output ports
	output [31:0] P;
	
	// Internal signals
	
	
endmodule
