`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// Create Date:    15:18:29 09/07/2012
// Module Name:    FBAddSub_LNCModule 
// Project Name: 	 Floating Point Project
// Author:			 Fredrik Brosser
//
// Description:	 Leading Nought Counter - Module for counting the number of leading
//						 noughts in a bit vector, i.e. #bits until first 1, starting from MSB
//
//////////////////////////////////////////////////////////////////////////////////

module FPAddSub_Pipelined_Simplified_2_0_LNCModule(
		A,
		Z
    );

	// Input ports
	input [25:0] A ;				// 32-bit input bit vector
	
	// Output ports
	output [4:0] Z ;				// Outputs number of leading noughts
	
	//reg [4:0] Z ;					// Outputs number of leading noughts
	wire [4:0] Z_in ;
	wire [15:0] val16 ;
	wire [7:0] val8 ;
	wire [3:0] val4 ;
	
	// Mapping to number of leading noughts (Ugly way to do this)
	/*
	assign Z_in[4] = (A[25:16] == 16'b0);
	assign val16     = Z_in[4] ? A[15:0] : A[25:16];
	assign Z_in[3] = (val16[15:8] == 8'b0);
	assign val8      = Z_in[3] ? val16[7:0] : val16[15:8];
	assign Z_in[2] = (val8[7:4] == 4'b0);
	assign val4      = Z_in[2] ? val8[3:0] : val8[7:4];
	assign Z_in[1] = (val4[3:2] == 2'b0);
	assign Z_in[0] = Z_in[1] ? ~val4[1] : ~val4[3];
	assign Z = Z_in ;
	*/
	/*
	assign Z = ( 
		A[25] ? 5'b00000 :	 
		A[24] ? 5'b00001 : 
		A[23] ? 5'b00010 : 
		A[22] ? 5'b00011 : 
		A[21] ? 5'b00100 : 
		A[20] ? 5'b00101 : 
		A[19] ? 5'b00110 : 
		A[18] ? 5'b00111 :
		A[17] ? 5'b01000 :
		A[16] ? 5'b01000 :
		A[15] ? 5'b01010 :
		A[14] ? 5'b01011 :
		A[13] ? 5'b01100 :
		A[12] ? 5'b01101 :
		A[11] ? 5'b01110 :
		A[10] ? 5'b01111 :
		A[9] ? 5'b10000 :
		A[8] ? 5'b10001 :
		A[7] ? 5'b10010 :
		A[6] ? 5'b10011 :
		A[5] ? 5'b10100 :
		A[4] ? 5'b10101 :
		A[3] ? 5'b10110 :
		A[2] ? 5'b10111 :
		A[1] ? 5'b11000 :
		A[0] ? 5'b11001 : 5'b11010
	);
	*/
	assign Z = ( 
		A[25] ? 0 :	 
		A[24] ? 1 : 
		A[23] ? 2 : 
		A[22] ? 3 : 
		A[21] ? 4 : 
		A[20] ? 5 : 
		A[19] ? 6 : 
		A[18] ? 7 :
		A[17] ? 8 :
		A[16] ? 9 :
		A[15] ? 10 :
		A[14] ? 11 :
		A[13] ? 12 :
		A[12] ? 13 :
		A[11] ? 14 :
		A[10] ? 15 :
		A[9] ? 16 :
		A[8] ? 17 :
		A[7] ? 18 :
		A[6] ? 19 :
		A[5] ? 20 :
		A[4] ? 21 :
		A[3] ? 22 :
		A[2] ? 23 :
		A[1] ? 24 :
		A[0] ? 25 : 26
	);
	/*
	always @(A) begin
		casez(A[25:0])
			26'b0: Z <= 26;
			26'b1: Z <= 25;
			26'b1?: Z <= 24;
			26'b1??: Z <= 23;
			26'b1???: Z <= 22;
			26'b1????: Z <= 21;
			26'b1?????: Z <= 20;
			26'b1??????: Z <= 19;
			26'b1???????: Z <= 18;
			26'b1????????: Z <= 17;
			26'b1?????????: Z <= 16;
			26'b1??????????: Z <= 15;
			26'b1???????????: Z <= 14;
			26'b1????????????: Z <= 13;
			26'b1?????????????: Z <= 12;
			26'b1??????????????: Z <= 11;
			26'b1???????????????: Z <= 10;
			26'b1????????????????: Z <= 9;
			26'b1?????????????????: Z <= 8;
			26'b1??????????????????: Z <= 7;
			26'b1???????????????????: Z <= 6;
			26'b1????????????????????: Z <= 5;
			26'b1?????????????????????: Z <= 4;
			26'b1??????????????????????: Z <= 3;
			26'b1???????????????????????: Z <= 2;
			26'b1????????????????????????: Z <= 1;
			26'b1?????????????????????????: Z <= 0;
			default : Z <= 0;
		endcase	
	end
	
	
	casez(A[25:0])
		26'b0: Z <= 26;
		26'b1: Z <= 25;
		26'b1?: Z <= 24;
		26'b1??: Z <= 23;
		26'b1???: Z <= 22;
		26'b1????: Z <= 21;
		26'b1?????: Z <= 20;
		26'b1??????: Z <= 19;
		26'b1???????: Z <= 18;
		26'b1????????: Z <= 17;
		26'b1?????????: Z <= 16;
		26'b1??????????: Z <= 15;
		26'b1???????????: Z <= 14;
		26'b1????????????: Z <= 13;
		26'b1?????????????: Z <= 12;
		26'b1??????????????: Z <= 11;
		26'b1???????????????: Z <= 10;
		26'b1????????????????: Z <= 9;
		26'b1?????????????????: Z <= 8;
		26'b1??????????????????: Z <= 7;
		26'b1???????????????????: Z <= 6;
		26'b1????????????????????: Z <= 5;
		26'b1?????????????????????: Z <= 4;
		26'b1??????????????????????: Z <= 3;
		26'b1???????????????????????: Z <= 2;
		26'b1????????????????????????: Z <= 1;
		26'b1?????????????????????????: Z <= 0;
		default : Z <= 0;
	endcase
	*/
	
endmodule
