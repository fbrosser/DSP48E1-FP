`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:00:37 09/10/2012
// Design Name:   FPAddSub
// Module Name:   P:/VerilogTraining/FPAddSub_Fred/FPAddSub_tb.v
// Project Name:  FPAddSub_Fred
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: FPAddSub
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module FPAddSub_tb;

	// Inputs
	reg clk;
	reg rst;
	reg [31:0] A;
	reg [31:0] B;
	reg Ctrl ;

	// Outputs
	wire [31:0] Z;
	wire [4:0] Flags;
	
	integer i ;
			
	// Instantiate the Unit Under Test (UUT)
	FPAddSub uut (
		.clk(clk),
		.rst(rst),
		.A(A), 
		.B(B), 
		.Ctrl(Ctrl),
		.Z(Z),
		.Flags(Flags)
	);

	always begin
		#5 clk = ~clk;
	end

	initial begin
		// Initialize Inputs
		A = 0;
		B = 0;
		clk = 0;
		Ctrl = 0;
		rst = 0;

		// Wait 100 ns for global reset to finish
		#10 rst = 1;
		#10 rst = 0;
        
		// Add stimulus here
		// 1+1 = 2 = 01000000000000000000000000000000
		#10 A = 32'b0_01111111_00000000000000000000000; B = 32'b0_01111111_00000000000000000000000; Ctrl = 1'b0;
		// 3+1 = 4 = 01000000100000000000000000000000
		#10 A = 32'b0_10000000_10000000000000000000000; B = 32'b0_01111111_00000000000000000000000; Ctrl = 1'b0;
		// 3+3 = 6 = 01000000110000000000000000000000
		#10 A = 32'b0_10000000_10000000000000000000000; B = 32'b0_10000000_10000000000000000000000; Ctrl = 1'b0;
		// 3.5+1.75 = 5.25 = 01000000101010000000000000000000 
		#10 A = 32'b0_10000000_11000000000000000000000; B = 32'b0_01111111_11000000000000000000000; Ctrl = 1'b0;
		// 28.0 + 0.15 = 28.15 = 01000001111000010011001100110011
		#10 A = 32'b0_10000011_11000000000000000000000 ; B = 32'b0_01111100_00110011001100110011010 ; Ctrl = 1'b0;
		// - 315.0 + -36.2	51 = -351.251 = 11000011101011111010000000100001
		#10 A = 32'b11000011100111011000000000000000 ; B = 32'b11000010000100010000000100000110 ; Ctrl = 1'b0; 
		// 832.312 - 23.1 = 809.212 = 01000100010010100100110110010001
		#10 A = 32'b01000100010100000001001111111000 ; B = 32'b01000001101110001100110011001101 ; Ctrl = 1'b1; 
		// 0.19 + 0.005 = 0.195 = 00111110010001111010111000010100
		#10 A = 32'b00111110010000101000111101011100 ; B = 32'b00111011101000111101011100001010 ; Ctrl = 1'b0; 
		// 0.1 + 0 = 0.1 = 00111101110011001100110011001101
		#10 A = 32'b00111101110011001100110011001101 ; B = 32'b00000000000000000000000000000000 ; Ctrl = 1'b0;
		// 28.0 + 0.15 = 28.15 = 01000001111000010011001100110011
		#10 A = 32'b01000001111000000000000000000000 ; B = 32'b00111110000110011001100110011010 ; Ctrl = 1'b0; 
		// - 12 - -0.07 = -11.93 = 11000001001111101110000101001000
		#10 A = 32'b11000001010000000000000000000000 ; B = 32'b10111101100011110101110000101001 ; Ctrl = 1'b1; 
		#9 $display("Z[12]: %b\n", Z);
		// -1252214.12412 + -125124 = -1377338.1 = 11001001101010000010000111010001
		#1 A = 32'b1_10010011_00110001101101110110001; B = 32'b1_10001111_11101000110001000000000; Ctrl = 1'b0; 
		#9 $display("Z[13]: %b\n", Z);
		// 100 + 0.000008 = 100.00001 = 01000010110010000000000000000001
		#1 A = 32'b0_10000101_10010000000000000000000; B = 32'b0_01101110_00001100011011110111101; Ctrl = 1'b0;
		#9 $display("Z[14]: %b\n", Z);
		// 1000 + 0.000008 = 1000 = 01000100011110100000000000000000
		#1 A = 32'b0_01111111_00000000000000000000000; B = 32'b0_01101110_00001100011011110111101; Ctrl = 1'b0;
		#9 $display("Z[15]: %b\n", Z);
		// 23672347 - 23672347 = 0 = 00000000000000000000000000000000
		#1 A = 32'b0_10010111_01101001001101100001110; B = 32'b0_10010111_01101001001101100001110; Ctrl = 1'b1; 
		#9 $display("Z[16]: %b\n", Z);
		// 23672347 + 23672347 = 47344694 = 01001100001101001001101100001110
		#1 A = 32'b0_10010111_01101001001101100001110; B = 32'b0_10010111_01101001001101100001110; Ctrl = 1'b0;  
		#9 $display("Z[17]: %b\n", Z);
		// 1 - 1 = 0 = 01001100001101001001101100001110
		#1 A = 32'b0_01111111_00000000000000000000000; B = 32'b0_01111111_00000000000000000000000; Ctrl = 1'b1;
		#9 $display("Z[18]: %b\n", Z);
		
		for (i=19; i<=28; i=i+1) begin
			#10 $display("Z[%d]: %b\n", i, Z);
		end
		
		#1000;
		#10 $finish;
		
	end
      
endmodule
