`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// Create Date:    01:56:20 09/07/2012 
// Module Name:    FPAddSub
// Project Name: 	 Floating Point Project
// Author:			 Fredrik Brosser
//
// Description:	 Top Module for a 32-bit floating point adder/subtractor.
//						 Follows the IEEE754 Single Precision standard.
//						 Supports only the default rounding mode.
//
//	Inputs:
//				a (32 bits)			: Single precision IEEE754 floating point number
//				b (32 bits)			: Single precision IEEE754 floating point number
//				operation (1 bit)	: Single control bit. 0/Addition, 1/Subtraction
//
//
// Outputs:
//				result (32 bits)	: Result of the operation, in IEEE754 Single format
//				flags	 (5 bits)	: Flags indicating exceptions:
//											Bit 4: Overflow
//											Bit 3: Underflow
//											Bit 2: Divide by Zero
//											Bit 1: Invalid/NaN
//											Bit 0: Inexact
//
//////////////////////////////////////////////////////////////////////////////////

module FPAddSub(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);
	
	// Clock and reset
	input clk ;						// Clock signal
	input rst ;						// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;				// Input A, a 32-bit floating point number
	input [31:0] b ;				// Input B, a 32-bit floating point number
	input operation ;					// Control signal
	
	// Output ports
	output [31:0] result ;				// result of the operation
	output [4:0] flags ;			// Flags indicating exceptions according to IEEE754
	
	// Pipeline Registers
	//reg [64:0] pipe_0;			// Pipeline register Input->PreAlign
	reg [81:0] pipe_1;			// Pipeline register PreAlign->Align1
	reg [78:0] pipe_2;			// Pipeline register Align1->Align3
	reg [78:0] pipe_3;			// Pipeline register Align1->Align3
	reg [71:0] pipe_4;			// Pipeline register Align3->Execute
	reg [51:0] pipe_5;			// Pipeline register Execute->Normalize
	reg [56:0] pipe_6;			// Pipeline register Nomalize->NormalizeShift1
	reg [56:0] pipe_8;			// Pipeline register NormalizeShift2->NormalizeShift3
	reg [54:0] pipe_9;		// Pipeline register NormalizeShift3->Round
	reg [41:0] pipe_10;			// Pipeline register NormalizeShift3->Round
	reg [36:0] pipe_11;			// Pipeline register NormalizeShift3->Round
	
	// Internal wires between modules
	wire [31:0] Aout_0 ;										// A's sign
	wire [31:0] Bout_0 ;										// B's sign
	wire Opout_0 ;										// A's sign
	
	wire Sa_0 ;										// A's sign
	wire Sb_0 ;										// B's sign
	wire MaxAB_0 ;									// Indicates the larger of A and B(0/A, 1/B)
	wire [7:0] CExp_0 ;							// Common Exponent
	wire [4:0] Shift_0 ;							// Number of steps to smaller mantissa shift right (align)
	wire [24:0] Mmax_0 ;							// Larger mantissa
	wire [4:0] InputExc_0 ;						// Input numbers are exceptions
	wire [9:0] ShiftDet_0 ;
	wire [31:0] MminS_0 ;						// Smaller mantissa after 0/16 shift
	
	wire [31:0] MminS_1 ;						// Smaller mantissa after 0/16 shift
	
	wire [31:0] MminS_2 ;						// Smaller mantissa after 0/4/8/12 shift
	
	wire [24:0] Mmin_3 ;							// Smaller mantissa after 0/1/2/3 shift
	wire G_3 ;										//Guard bit
	wire PS_3 ;										// Pre-sticky bit
	
	wire [32:0] Sum_4 ;
	wire PSgn_4 ;
	wire Opr_4 ;
	
	wire [4:0] Shift_5 ;							// Number of steps to shift sum left (normalize)
	wire [32:0] SumS_5 ;							// Sum after 0/16 shift

	wire [32:0] SumS_6 ;							// Sum after 0/16 shift
	
	wire [32:0] SumS_7 ;							// Sum after 0/16 shift
	
	wire [22:0] NormM_8 ;							// Normalized mantissa
	wire [8:0] NormE_8;							// Adjusted exponent
	
	wire ZeroSum_8 ;								// Zero flag
	wire NegE_8 ;									// Flag indicating negative exponent
	wire R_8 ;										// Round bit
	wire S_8 ;										// Final sticky bit
	wire FG_8 ;										// Final sticky bit
	
	wire [31:0] P_int ;
	//wire [31:0] Z_int ;
	wire EOF ;
	//wire [4:0] Flags_int ;
	
	//assign result = pipe_11[31:0] ;
	//assign flags = pipe_11[36:32] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_PrealignModule PrealignModule
	(	
		// Inputs
		a, b, operation,
		//pipe_0[63:32], pipe_0[31:0],
		// Outputs
		Sa_0, Sb_0, ShiftDet_0[9:0], InputExc_0[4:0], Aout_0[31:0], Bout_0[31:0], Opout_0
	) ;
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_AlignModule AlignModule
	(	
		// Inputs
		pipe_1[80:49], pipe_1[48:17], pipe_1[14:5],
		// Outputs
		CExp_0[7:0], MaxAB_0, Shift_0[4:0], MminS_0[31:0], Mmax_0[24:0]
	) ;	
	// Alignment Shift Stage 1
	FPAddSub_AlignShift1 AlignShift1
	(
		// Inputs
		pipe_2[31:0], pipe_2[66:62],
		// Outputs
		MminS_2[31:0]                
	) ;

	// Alignment Shift Stage 3 and compution of guard and sticky bits
	FPAddSub_AlignShift2 AlignShift2
	(
		// Inputs
		pipe_3[31:0], pipe_3[66:62],
		// Outputs
		Mmin_3[24:0]
	) ;
	// Perform mantissa addition
	FPAddSub_ExecutionModule ExecutionModule
	(
		// Inputs
		pipe_4[54:30], pipe_4[24:0], pipe_4[70], pipe_4[69], pipe_4[68], pipe_4[71],
		// Outputs
		Sum_4[32:0], PSgn_4, Opr_4
	) ;
	
	// Prepare normalization of result
	FPAddSub_NormalizeModule NormalizeModule
	(
		// Inputs
		pipe_5[32:0], 
		// Outputs
		SumS_5[32:0], Shift_5[4:0]
		) ;
					
	// Normalization Shift Stage 1
	FPAddSub_NormalizeShift1 NormalizeShift1
	(
		// Inputs
		pipe_6[32:0], pipe_6[55:51],
		// Outputs
		SumS_7[32:0]
	) ;
		
	// Normalization Shift Stage 3 and final guard, sticky and round bits
	FPAddSub_NormalizeShift2 NormalizeShift2
	(
		// Inputs
		pipe_8[32:0],
		pipe_8[45:38],
		pipe_8[49],
		pipe_8[55:51],
		// Outputs
		NormM_8[22:0],					// Normalized mantissa
		NormE_8[8:0],					// Adjusted exponent
		ZeroSum_8,						// Zero flag
		NegE_8,							// Flag indicating negative exponent
		R_8,								// Round bit
		S_8,								// Final sticky bit
		FG_8
	) ;

	// Round and put result together
	FPAddSub_RoundModule RoundModule
	(
		// Inputs
		 pipe_9[3], pipe_9[52], pipe_9[12:4], pipe_9[35:13], pipe_9[1], pipe_9[0], pipe_9[54], pipe_9[51], pipe_9[50], pipe_9[53], pipe_9[49], 
		// Outputs
		P_int[31:0], EOF
	) ;
	
	// Check for exceptions
	FPAddSub_ExceptionModule Exceptionmodule
	(
		// Inputs
		pipe_10[40:9], pipe_10[41], pipe_10[8], pipe_10[7], pipe_10[6], pipe_10[5:1], pipe_10[0], 
		// Outputs
		result[31:0],
		flags[4:0]
		//Z_int[31:0],
		//Flags_int[4:0]
	) ;			
	
	always @ (posedge clk) begin	
		if(rst) begin
			//pipe_0 <= 0;
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
			pipe_4 <= 0;
			pipe_5 <= 0;
			pipe_6 <= 0;
			pipe_8 <= 0;
			pipe_9 <= 0;
			pipe_10 <= 0;
		end 
		else begin
		
			/* PIPE_0 :
				[64] operation
				[63:32] A
				[31:0] B
			*/
			//pipe_0 <= {operation, a, b} ;	
			/* PIPE_1 :
				[81] operation
				[80:49] A
				[48:17] B
				[16] Sa_0
				[15] Sb_0
				[14:5] ShiftDet
				[4:0] InputExc_0
			*/
			pipe_1 <= {Opout_0, Aout_0[31:0], Bout_0[31:0], Sa_0, Sb_0, ShiftDet_0[9:0], InputExc_0[4:0]} ;	
			/* PIPE_2 :
				[78] operation
				[77] Sa_0
				[76] Sb_0
				[75] MaxAB_0
				[74:67] CExp_0
				[66:62] Shift_0
				[61:37] Mmax_0
				[36:32] InputExc_0
				[31:0] MminS_1
			*/
			pipe_2 <= {pipe_1[81], pipe_1[16:15], MaxAB_0, CExp_0[7:0], Shift_0[4:0], Mmax_0[24:0], pipe_1[4:0], MminS_0[31:0]} ;	
			/* PIPE_3 :
				[78] operation
				[77] Sa_0
				[76] Sb_0
				[75] MaxAB_0
				[74:67] CExp_0
				[66:62] Shift_0
				[61:37] Mmax_0
				[36:32] InputExc_0
				[31:0] MminS_1
			*/
			pipe_3 <= {pipe_2[78:32], MminS_2[31:0]} ;	
			/* PIPE_4 :
				[71] operation
				[70] Sa_0
				[69] Sb_0
				[68] MaxAB_0
				[67:60] CExp_0
				[59:55] Shift_0
				[54:30] Mmax_0
				[29:25] InputExc_0
				[24:0] Mmin_3
			*/					
			pipe_4 <= {pipe_3[78:32], Mmin_3[24:0]} ;	
			/* PIPE_5 :
				[51] operation
				[50] PSgn_4
				[49] Opr_4
				[48] Sa_0
				[47] Sb_0
				[46] MaxAB_0
				[45:38] CExp_0
				[37:33] InputExc_0
				[32:0] Sum_4
			*/					
			pipe_5 <= {pipe_4[71], PSgn_4, Opr_4, pipe_4[70:60], pipe_4[29:25], Sum_4[32:0]} ;
			/* PIPE_6 :
				[56] operation
				[55:51] Shift_5
				[50] PSgn_4
				[49] Opr_4
				[48] Sa_0
				[47] Sb_0
				[46] MaxAB_0
				[45:38] CExp_0
				[37:33] InputExc_0
				[32:0] Sum_4
			*/					
			pipe_6 <= {pipe_5[51], Shift_5[4:0], pipe_5[50:33], SumS_5[32:0]} ;	
			/* PIPE_8 :
				[56] operation
				[55:51] Shift_5
				[50] PSgn_4
				[49] Opr_4
				[48] Sa_0
				[47] Sb_0
				[46] MaxAB_0
				[45:38] CExp_0
				[37:33] InputExc_0
				[32:0] Sum_4
			*/						
			pipe_8 <= {pipe_6[56:33], SumS_7[32:0]} ;	
			/* PIPE_9:
				[54] FG_8 
				[53] operation
				[52] PSgn_4
				[51] Sa_0
				[50] Sb_0
				[49] MaxAB_0
				[48:41] CExp_0
				[40:36] InputExc_8
				[35:13] NormM_8 
				[12:4] NormE_8
				[3] ZeroSum_8
				[2] NegE_8
				[1] R_8
				[0] S_8
			*/				
			pipe_9 <= {FG_8, pipe_8[56], pipe_8[50], pipe_8[48:33], NormM_8[22:0], NormE_8[8:0], ZeroSum_8, NegE_8, R_8, S_8} ;	
			/* PIPE_10:
				[41] ZeroSum
				[40:9] P_int
				[8] NegE_8
				[7] R_8
				[6] S_8
				[5:1] InputExc_8
				[0] EOF
			*/				
			pipe_10 <= {pipe_9[3], P_int[31:0], pipe_9[2], pipe_9[1], pipe_9[0], pipe_9[40:36], EOF} ;	
			/*
				PIPE_11:
				[36:32] Flags
				[31:0]  result
			*/
			//pipe_11 <= {Flags_int[4:0], Z_int[31:0]} ;	
		end
	end		

endmodule
