`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   23:24:54 09/20/2012
// Design Name:   FPMult
// Module Name:   P:/VerilogTraining/FPMult/FPMult_tb.v
// Project Name:  FPMult
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: FPMult
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module FPMult_tb;

	// Inputs
	reg [31:0] A;
	reg [31:0] B;
	reg [2:0] Ctrl;

	// Outputs
	wire [31:0] P;

	// Instantiate the Unit Under Test (UUT)
	FPMult uut (
		.A(A), 
		.B(B), 
		.Ctrl(Ctrl),
		.P(P)
	);

	initial begin
		// Initialize Inputs
		A = 0;
		B = 0;
		Ctrl = 0;

		// Wait 100 ns for global reset to finish
		#10;
        
		// Add stimulus here
		// 2.5 * 4.75 = 11.875 = 		01000001001111100000000000000000
		#10 A = 32'b0__1000_0000__0100_0000_0000_0000_0000_000; B = 32'b0__1000_0001__0011_0000_0000_0000_0000_000;
		#10 $display("P[1]: %b\n", P);
		
		// 1 * 1 = 1 = 					00111111100000000000000000000000
		//										00111111100000000000000000000000
		#10 A = 32'b0__0111_1111__0000_0000_0000_0000_0000_000; B = 32'b0__0111_1111__0000_0000_0000_0000_0000_000;
		#10 $display("P[2]: %b\n", P);
		
		// 3 * 2 = 6 = 					01000000110000000000000000000000
		//										01000000110000000000000000000000
		#10 A = 32'b0__1000_0000__1000_0000_0000_0000_0000_000; B = 32'b0__1000_0000__0000_0000_0000_0000_0000_000;
		#10 $display("P[3]: %b\n", P);
		
		// 2 * -3 = -6 = 					11000000110000000000000000000000
		//										11000000110000000000000000000000
		#10 A = 32'b0__1000_0000__1000_0000_0000_0000_0000_000; B = 32'b1__1000_0000__0000_0000_0000_0000_0000_000;
		#10 $display("P[4]: %b\n", P);
		
		// 14.56 * -23.1351 = -336.84705 = 	11000011101010000110110001101100
		//												11000011101010000110110001101100
		#10 A = 32'b01000001011010001111010111000011; B = 32'b11000001101110010001010010101111;
		#10 $display("P[5]: %b\n", P);
		
		// - 12 * -0.07 = 0.84 = 		00111111010101110000101000111101
		//										00111111010101110000101000111110
		#10 A = 32'b11000001010000000000000000000000 ; B = 32'b10111101100011110101110000101001 ; 
		#10 $display("P[6]: %b\n", P);
		
		// - 315.0 * -36.251 = 11419.065 = 	01000110001100100110110001000011
		//												01000110001100100110110001000010
		#10 A = 32'b11000011100111011000000000000000 ; B = 32'b11000010000100010000000100000110 ;
		#10 $display("P[7]: %b\n", P);
		
		// 832.312 * 23.1 = 19226.4072 = 	01000110100101100011010011010000
		//												01000110100101100011010011010001
		#10 A = 32'b01000100010100000001001111111000 ; B = 32'b01000001101110001100110011001101 ; 
		#10 $display("P[8]: %b\n", P);
		
		#10 $finish;
	end
      
endmodule

